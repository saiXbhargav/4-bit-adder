magic
tech scmos
timestamp 1731995772
<< nwell >>
rect 517 -474 541 -450
rect 556 -460 590 -454
rect 657 -457 681 -433
rect 696 -443 730 -437
rect 556 -490 618 -460
rect 696 -473 758 -443
rect 792 -457 816 -433
rect 831 -443 865 -437
rect 831 -473 893 -443
rect 930 -458 954 -434
rect 969 -444 1003 -438
rect 724 -479 758 -473
rect 859 -479 893 -473
rect 969 -474 1031 -444
rect 997 -480 1031 -474
rect 584 -496 618 -490
rect 517 -529 541 -505
rect 657 -512 681 -488
rect 792 -512 816 -488
rect 930 -513 954 -489
rect 442 -601 479 -575
rect 485 -601 513 -575
rect 649 -588 677 -562
rect 685 -587 713 -561
rect 723 -587 751 -561
rect 762 -588 790 -562
rect 811 -594 839 -568
rect 879 -601 903 -577
rect 918 -587 952 -581
rect 918 -617 980 -587
rect 946 -623 980 -617
rect 442 -675 479 -649
rect 485 -675 513 -649
rect 816 -670 844 -644
rect 879 -656 903 -632
rect 442 -744 479 -718
rect 485 -744 513 -718
rect 819 -746 847 -720
rect 890 -737 914 -713
rect 929 -723 963 -717
rect 929 -753 991 -723
rect 957 -759 991 -753
rect 890 -792 914 -768
rect 442 -818 479 -792
rect 485 -818 513 -792
rect 820 -818 848 -792
rect 899 -871 923 -847
rect 938 -857 972 -851
rect 479 -904 507 -878
rect 938 -887 1000 -857
rect 966 -893 1000 -887
rect 899 -926 923 -902
rect 904 -1020 928 -996
rect 943 -1006 977 -1000
rect 943 -1036 1005 -1006
rect 971 -1042 1005 -1036
rect 904 -1075 928 -1051
<< ntransistor >>
rect 528 -488 530 -482
rect 668 -471 670 -465
rect 803 -471 805 -465
rect 941 -472 943 -466
rect 707 -520 709 -508
rect 717 -520 719 -508
rect 735 -520 737 -508
rect 745 -520 747 -508
rect 842 -520 844 -508
rect 852 -520 854 -508
rect 870 -520 872 -508
rect 880 -520 882 -508
rect 567 -537 569 -525
rect 577 -537 579 -525
rect 595 -537 597 -525
rect 605 -537 607 -525
rect 668 -526 670 -520
rect 803 -526 805 -520
rect 980 -521 982 -509
rect 990 -521 992 -509
rect 1008 -521 1010 -509
rect 1018 -521 1020 -509
rect 941 -527 943 -521
rect 528 -543 530 -537
rect 823 -611 825 -604
rect 455 -629 457 -616
rect 465 -629 467 -616
rect 497 -618 499 -611
rect 890 -615 892 -609
rect 455 -703 457 -690
rect 465 -703 467 -690
rect 497 -692 499 -685
rect 455 -772 457 -759
rect 465 -772 467 -759
rect 497 -761 499 -754
rect 455 -846 457 -833
rect 465 -846 467 -833
rect 497 -835 499 -828
rect 553 -836 555 -623
rect 560 -836 562 -623
rect 607 -835 609 -622
rect 640 -835 642 -622
rect 671 -835 673 -622
rect 705 -834 707 -621
rect 726 -834 728 -621
rect 748 -834 750 -621
rect 776 -833 778 -620
rect 929 -664 931 -652
rect 939 -664 941 -652
rect 957 -664 959 -652
rect 967 -664 969 -652
rect 890 -670 892 -664
rect 828 -687 830 -680
rect 901 -751 903 -745
rect 831 -763 833 -756
rect 940 -800 942 -788
rect 950 -800 952 -788
rect 968 -800 970 -788
rect 978 -800 980 -788
rect 901 -806 903 -800
rect 832 -835 834 -828
rect 910 -885 912 -879
rect 491 -921 493 -914
rect 949 -934 951 -922
rect 959 -934 961 -922
rect 977 -934 979 -922
rect 987 -934 989 -922
rect 910 -940 912 -934
rect 344 -973 548 -971
rect 915 -1034 917 -1028
rect 954 -1083 956 -1071
rect 964 -1083 966 -1071
rect 982 -1083 984 -1071
rect 992 -1083 994 -1071
rect 915 -1089 917 -1083
<< ptransistor >>
rect 668 -451 670 -439
rect 528 -468 530 -456
rect 567 -484 569 -460
rect 577 -484 579 -460
rect 595 -490 597 -466
rect 605 -490 607 -466
rect 707 -467 709 -443
rect 717 -467 719 -443
rect 735 -473 737 -449
rect 745 -473 747 -449
rect 803 -451 805 -439
rect 842 -467 844 -443
rect 852 -467 854 -443
rect 528 -523 530 -511
rect 668 -506 670 -494
rect 870 -473 872 -449
rect 880 -473 882 -449
rect 941 -452 943 -440
rect 980 -468 982 -444
rect 990 -468 992 -444
rect 803 -506 805 -494
rect 1008 -474 1010 -450
rect 1018 -474 1020 -450
rect 941 -507 943 -495
rect 661 -580 663 -568
rect 697 -579 699 -567
rect 735 -579 737 -567
rect 455 -593 457 -581
rect 465 -593 467 -581
rect 497 -593 499 -581
rect 774 -580 776 -568
rect 823 -586 825 -574
rect 890 -595 892 -583
rect 929 -611 931 -587
rect 939 -611 941 -587
rect 455 -667 457 -655
rect 465 -667 467 -655
rect 497 -667 499 -655
rect 455 -736 457 -724
rect 465 -736 467 -724
rect 497 -736 499 -724
rect 455 -810 457 -798
rect 465 -810 467 -798
rect 497 -810 499 -798
rect 957 -617 959 -593
rect 967 -617 969 -593
rect 890 -650 892 -638
rect 828 -662 830 -650
rect 831 -738 833 -726
rect 901 -731 903 -719
rect 940 -747 942 -723
rect 950 -747 952 -723
rect 968 -753 970 -729
rect 978 -753 980 -729
rect 901 -786 903 -774
rect 832 -810 834 -798
rect 910 -865 912 -853
rect 491 -896 493 -884
rect 949 -881 951 -857
rect 959 -881 961 -857
rect 977 -887 979 -863
rect 987 -887 989 -863
rect 910 -920 912 -908
rect 915 -1014 917 -1002
rect 954 -1030 956 -1006
rect 964 -1030 966 -1006
rect 982 -1036 984 -1012
rect 992 -1036 994 -1012
rect 915 -1069 917 -1057
<< ndiffusion >>
rect 527 -488 528 -482
rect 530 -488 531 -482
rect 667 -471 668 -465
rect 670 -471 671 -465
rect 802 -471 803 -465
rect 805 -471 806 -465
rect 940 -472 941 -466
rect 943 -472 944 -466
rect 706 -520 707 -508
rect 709 -520 717 -508
rect 719 -520 720 -508
rect 734 -520 735 -508
rect 737 -520 745 -508
rect 747 -520 748 -508
rect 841 -520 842 -508
rect 844 -520 852 -508
rect 854 -520 855 -508
rect 869 -520 870 -508
rect 872 -520 880 -508
rect 882 -520 883 -508
rect 566 -537 567 -525
rect 569 -537 577 -525
rect 579 -537 580 -525
rect 594 -537 595 -525
rect 597 -537 605 -525
rect 607 -537 608 -525
rect 667 -526 668 -520
rect 670 -526 671 -520
rect 802 -526 803 -520
rect 805 -526 806 -520
rect 979 -521 980 -509
rect 982 -521 990 -509
rect 992 -521 993 -509
rect 1007 -521 1008 -509
rect 1010 -521 1018 -509
rect 1020 -521 1021 -509
rect 940 -527 941 -521
rect 943 -527 944 -521
rect 527 -543 528 -537
rect 530 -543 531 -537
rect 822 -611 823 -604
rect 825 -611 826 -604
rect 454 -629 455 -616
rect 457 -629 465 -616
rect 467 -629 468 -616
rect 496 -618 497 -611
rect 499 -618 500 -611
rect 889 -615 890 -609
rect 892 -615 893 -609
rect 454 -703 455 -690
rect 457 -703 465 -690
rect 467 -703 468 -690
rect 496 -692 497 -685
rect 499 -692 500 -685
rect 454 -772 455 -759
rect 457 -772 465 -759
rect 467 -772 468 -759
rect 496 -761 497 -754
rect 499 -761 500 -754
rect 454 -846 455 -833
rect 457 -846 465 -833
rect 467 -846 468 -833
rect 496 -835 497 -828
rect 499 -835 500 -828
rect 552 -836 553 -623
rect 555 -836 560 -623
rect 562 -836 563 -623
rect 606 -835 607 -622
rect 609 -835 610 -622
rect 639 -835 640 -622
rect 642 -835 643 -622
rect 670 -835 671 -622
rect 673 -835 674 -622
rect 704 -834 705 -621
rect 707 -834 708 -621
rect 725 -834 726 -621
rect 728 -834 729 -621
rect 747 -834 748 -621
rect 750 -834 751 -621
rect 775 -833 776 -620
rect 778 -833 779 -620
rect 928 -664 929 -652
rect 931 -664 939 -652
rect 941 -664 942 -652
rect 956 -664 957 -652
rect 959 -664 967 -652
rect 969 -664 970 -652
rect 889 -670 890 -664
rect 892 -670 893 -664
rect 827 -687 828 -680
rect 830 -687 831 -680
rect 900 -751 901 -745
rect 903 -751 904 -745
rect 830 -763 831 -756
rect 833 -763 834 -756
rect 939 -800 940 -788
rect 942 -800 950 -788
rect 952 -800 953 -788
rect 967 -800 968 -788
rect 970 -800 978 -788
rect 980 -800 981 -788
rect 900 -806 901 -800
rect 903 -806 904 -800
rect 831 -835 832 -828
rect 834 -835 835 -828
rect 909 -885 910 -879
rect 912 -885 913 -879
rect 490 -921 491 -914
rect 493 -921 494 -914
rect 948 -934 949 -922
rect 951 -934 959 -922
rect 961 -934 962 -922
rect 976 -934 977 -922
rect 979 -934 987 -922
rect 989 -934 990 -922
rect 909 -940 910 -934
rect 912 -940 913 -934
rect 344 -971 548 -970
rect 344 -974 548 -973
rect 914 -1034 915 -1028
rect 917 -1034 918 -1028
rect 953 -1083 954 -1071
rect 956 -1083 964 -1071
rect 966 -1083 967 -1071
rect 981 -1083 982 -1071
rect 984 -1083 992 -1071
rect 994 -1083 995 -1071
rect 914 -1089 915 -1083
rect 917 -1089 918 -1083
<< pdiffusion >>
rect 667 -451 668 -439
rect 670 -451 671 -439
rect 527 -468 528 -456
rect 530 -468 531 -456
rect 566 -484 567 -460
rect 569 -484 571 -460
rect 575 -484 577 -460
rect 579 -484 580 -460
rect 594 -490 595 -466
rect 597 -490 599 -466
rect 603 -490 605 -466
rect 607 -490 608 -466
rect 706 -467 707 -443
rect 709 -467 711 -443
rect 715 -467 717 -443
rect 719 -467 720 -443
rect 734 -473 735 -449
rect 737 -473 739 -449
rect 743 -473 745 -449
rect 747 -473 748 -449
rect 802 -451 803 -439
rect 805 -451 806 -439
rect 841 -467 842 -443
rect 844 -467 846 -443
rect 850 -467 852 -443
rect 854 -467 855 -443
rect 527 -523 528 -511
rect 530 -523 531 -511
rect 667 -506 668 -494
rect 670 -506 671 -494
rect 869 -473 870 -449
rect 872 -473 874 -449
rect 878 -473 880 -449
rect 882 -473 883 -449
rect 940 -452 941 -440
rect 943 -452 944 -440
rect 979 -468 980 -444
rect 982 -468 984 -444
rect 988 -468 990 -444
rect 992 -468 993 -444
rect 802 -506 803 -494
rect 805 -506 806 -494
rect 1007 -474 1008 -450
rect 1010 -474 1012 -450
rect 1016 -474 1018 -450
rect 1020 -474 1021 -450
rect 940 -507 941 -495
rect 943 -507 944 -495
rect 660 -580 661 -568
rect 663 -580 664 -568
rect 696 -579 697 -567
rect 699 -579 700 -567
rect 734 -579 735 -567
rect 737 -579 738 -567
rect 454 -593 455 -581
rect 457 -593 459 -581
rect 463 -593 465 -581
rect 467 -593 468 -581
rect 496 -593 497 -581
rect 499 -593 500 -581
rect 773 -580 774 -568
rect 776 -580 777 -568
rect 822 -586 823 -574
rect 825 -586 826 -574
rect 889 -595 890 -583
rect 892 -595 893 -583
rect 928 -611 929 -587
rect 931 -611 933 -587
rect 937 -611 939 -587
rect 941 -611 942 -587
rect 454 -667 455 -655
rect 457 -667 459 -655
rect 463 -667 465 -655
rect 467 -667 468 -655
rect 496 -667 497 -655
rect 499 -667 500 -655
rect 454 -736 455 -724
rect 457 -736 459 -724
rect 463 -736 465 -724
rect 467 -736 468 -724
rect 496 -736 497 -724
rect 499 -736 500 -724
rect 454 -810 455 -798
rect 457 -810 459 -798
rect 463 -810 465 -798
rect 467 -810 468 -798
rect 496 -810 497 -798
rect 499 -810 500 -798
rect 956 -617 957 -593
rect 959 -617 961 -593
rect 965 -617 967 -593
rect 969 -617 970 -593
rect 889 -650 890 -638
rect 892 -650 893 -638
rect 827 -662 828 -650
rect 830 -662 831 -650
rect 830 -738 831 -726
rect 833 -738 834 -726
rect 900 -731 901 -719
rect 903 -731 904 -719
rect 939 -747 940 -723
rect 942 -747 944 -723
rect 948 -747 950 -723
rect 952 -747 953 -723
rect 967 -753 968 -729
rect 970 -753 972 -729
rect 976 -753 978 -729
rect 980 -753 981 -729
rect 900 -786 901 -774
rect 903 -786 904 -774
rect 831 -810 832 -798
rect 834 -810 835 -798
rect 909 -865 910 -853
rect 912 -865 913 -853
rect 490 -896 491 -884
rect 493 -896 494 -884
rect 948 -881 949 -857
rect 951 -881 953 -857
rect 957 -881 959 -857
rect 961 -881 962 -857
rect 976 -887 977 -863
rect 979 -887 981 -863
rect 985 -887 987 -863
rect 989 -887 990 -863
rect 909 -920 910 -908
rect 912 -920 913 -908
rect 914 -1014 915 -1002
rect 917 -1014 918 -1002
rect 953 -1030 954 -1006
rect 956 -1030 958 -1006
rect 962 -1030 964 -1006
rect 966 -1030 967 -1006
rect 981 -1036 982 -1012
rect 984 -1036 986 -1012
rect 990 -1036 992 -1012
rect 994 -1036 995 -1012
rect 914 -1069 915 -1057
rect 917 -1069 918 -1057
<< ndcontact >>
rect 523 -488 527 -482
rect 531 -488 535 -482
rect 663 -471 667 -465
rect 671 -471 675 -465
rect 798 -471 802 -465
rect 806 -471 810 -465
rect 936 -472 940 -466
rect 944 -472 948 -466
rect 702 -520 706 -508
rect 720 -520 724 -508
rect 730 -520 734 -508
rect 748 -520 752 -508
rect 837 -520 841 -508
rect 855 -520 859 -508
rect 865 -520 869 -508
rect 883 -520 887 -508
rect 562 -537 566 -525
rect 580 -537 584 -525
rect 590 -537 594 -525
rect 608 -537 612 -525
rect 663 -526 667 -520
rect 671 -526 675 -520
rect 798 -526 802 -520
rect 806 -526 810 -520
rect 975 -521 979 -509
rect 993 -521 997 -509
rect 1003 -521 1007 -509
rect 1021 -521 1025 -509
rect 936 -527 940 -521
rect 944 -527 948 -521
rect 523 -543 527 -537
rect 531 -543 535 -537
rect 818 -611 822 -604
rect 826 -611 830 -604
rect 450 -629 454 -616
rect 468 -629 472 -616
rect 492 -618 496 -611
rect 500 -618 504 -611
rect 885 -615 889 -609
rect 893 -615 897 -609
rect 450 -703 454 -690
rect 468 -703 472 -690
rect 492 -692 496 -685
rect 500 -692 504 -685
rect 450 -772 454 -759
rect 468 -772 472 -759
rect 492 -761 496 -754
rect 500 -761 504 -754
rect 450 -846 454 -833
rect 468 -846 472 -833
rect 492 -835 496 -828
rect 500 -835 504 -828
rect 548 -836 552 -623
rect 563 -836 568 -623
rect 602 -835 606 -622
rect 610 -835 614 -622
rect 635 -835 639 -622
rect 643 -835 647 -622
rect 666 -835 670 -622
rect 674 -835 678 -622
rect 700 -834 704 -621
rect 708 -834 712 -621
rect 721 -834 725 -621
rect 729 -834 733 -621
rect 743 -834 747 -621
rect 751 -834 755 -621
rect 771 -833 775 -620
rect 779 -833 783 -620
rect 924 -664 928 -652
rect 942 -664 946 -652
rect 952 -664 956 -652
rect 970 -664 974 -652
rect 885 -670 889 -664
rect 893 -670 897 -664
rect 823 -687 827 -680
rect 831 -687 835 -680
rect 896 -751 900 -745
rect 904 -751 908 -745
rect 826 -763 830 -756
rect 834 -763 838 -756
rect 935 -800 939 -788
rect 953 -800 957 -788
rect 963 -800 967 -788
rect 981 -800 985 -788
rect 896 -806 900 -800
rect 904 -806 908 -800
rect 827 -835 831 -828
rect 835 -835 839 -828
rect 905 -885 909 -879
rect 913 -885 917 -879
rect 486 -921 490 -914
rect 494 -921 498 -914
rect 944 -934 948 -922
rect 962 -934 966 -922
rect 972 -934 976 -922
rect 990 -934 994 -922
rect 905 -940 909 -934
rect 913 -940 917 -934
rect 344 -970 548 -966
rect 344 -978 548 -974
rect 910 -1034 914 -1028
rect 918 -1034 922 -1028
rect 949 -1083 953 -1071
rect 967 -1083 971 -1071
rect 977 -1083 981 -1071
rect 995 -1083 999 -1071
rect 910 -1089 914 -1083
rect 918 -1089 922 -1083
<< pdcontact >>
rect 663 -451 667 -439
rect 671 -451 675 -439
rect 523 -468 527 -456
rect 531 -468 535 -456
rect 562 -484 566 -460
rect 571 -484 575 -460
rect 580 -484 584 -460
rect 590 -490 594 -466
rect 599 -490 603 -466
rect 608 -490 612 -466
rect 702 -467 706 -443
rect 711 -467 715 -443
rect 720 -467 724 -443
rect 730 -473 734 -449
rect 739 -473 743 -449
rect 748 -473 752 -449
rect 798 -451 802 -439
rect 806 -451 810 -439
rect 837 -467 841 -443
rect 846 -467 850 -443
rect 855 -467 859 -443
rect 523 -523 527 -511
rect 531 -523 535 -511
rect 663 -506 667 -494
rect 671 -506 675 -494
rect 865 -473 869 -449
rect 874 -473 878 -449
rect 883 -473 887 -449
rect 936 -452 940 -440
rect 944 -452 948 -440
rect 975 -468 979 -444
rect 984 -468 988 -444
rect 993 -468 997 -444
rect 798 -506 802 -494
rect 806 -506 810 -494
rect 1003 -474 1007 -450
rect 1012 -474 1016 -450
rect 1021 -474 1025 -450
rect 936 -507 940 -495
rect 944 -507 948 -495
rect 656 -580 660 -568
rect 664 -580 668 -568
rect 692 -579 696 -567
rect 700 -579 704 -567
rect 730 -579 734 -567
rect 738 -579 742 -567
rect 450 -593 454 -581
rect 459 -593 463 -581
rect 468 -593 472 -581
rect 492 -593 496 -581
rect 500 -593 504 -581
rect 769 -580 773 -568
rect 777 -580 781 -568
rect 818 -586 822 -574
rect 826 -586 830 -574
rect 885 -595 889 -583
rect 893 -595 897 -583
rect 924 -611 928 -587
rect 933 -611 937 -587
rect 942 -611 946 -587
rect 450 -667 454 -655
rect 459 -667 463 -655
rect 468 -667 472 -655
rect 492 -667 496 -655
rect 500 -667 504 -655
rect 450 -736 454 -724
rect 459 -736 463 -724
rect 468 -736 472 -724
rect 492 -736 496 -724
rect 500 -736 504 -724
rect 450 -810 454 -798
rect 459 -810 463 -798
rect 468 -810 472 -798
rect 492 -810 496 -798
rect 500 -810 504 -798
rect 952 -617 956 -593
rect 961 -617 965 -593
rect 970 -617 974 -593
rect 885 -650 889 -638
rect 893 -650 897 -638
rect 823 -662 827 -650
rect 831 -662 835 -650
rect 826 -738 830 -726
rect 834 -738 838 -726
rect 896 -731 900 -719
rect 904 -731 908 -719
rect 935 -747 939 -723
rect 944 -747 948 -723
rect 953 -747 957 -723
rect 963 -753 967 -729
rect 972 -753 976 -729
rect 981 -753 985 -729
rect 896 -786 900 -774
rect 904 -786 908 -774
rect 827 -810 831 -798
rect 835 -810 839 -798
rect 905 -865 909 -853
rect 913 -865 917 -853
rect 486 -896 490 -884
rect 494 -896 498 -884
rect 944 -881 948 -857
rect 953 -881 957 -857
rect 962 -881 966 -857
rect 972 -887 976 -863
rect 981 -887 985 -863
rect 990 -887 994 -863
rect 905 -920 909 -908
rect 913 -920 917 -908
rect 910 -1014 914 -1002
rect 918 -1014 922 -1002
rect 949 -1030 953 -1006
rect 958 -1030 962 -1006
rect 967 -1030 971 -1006
rect 977 -1036 981 -1012
rect 986 -1036 990 -1012
rect 995 -1036 999 -1012
rect 910 -1069 914 -1057
rect 918 -1069 922 -1057
<< polysilicon >>
rect 668 -439 670 -436
rect 803 -439 805 -436
rect 707 -443 709 -440
rect 717 -443 719 -440
rect 528 -456 530 -453
rect 567 -460 569 -457
rect 577 -460 579 -457
rect 528 -482 530 -468
rect 595 -466 597 -463
rect 605 -466 607 -463
rect 668 -465 670 -451
rect 528 -491 530 -488
rect 567 -493 569 -484
rect 577 -494 579 -484
rect 735 -449 737 -446
rect 745 -449 747 -446
rect 668 -474 670 -471
rect 707 -476 709 -467
rect 717 -477 719 -467
rect 941 -440 943 -437
rect 842 -443 844 -440
rect 852 -443 854 -440
rect 803 -465 805 -451
rect 870 -449 872 -446
rect 880 -449 882 -446
rect 528 -511 530 -508
rect 528 -537 530 -523
rect 567 -525 569 -498
rect 577 -525 579 -499
rect 595 -501 597 -490
rect 595 -525 597 -505
rect 605 -512 607 -490
rect 668 -494 670 -491
rect 605 -525 607 -516
rect 668 -520 670 -506
rect 707 -508 709 -481
rect 717 -508 719 -482
rect 735 -484 737 -473
rect 735 -508 737 -488
rect 745 -495 747 -473
rect 803 -474 805 -471
rect 842 -476 844 -467
rect 852 -477 854 -467
rect 980 -444 982 -441
rect 990 -444 992 -441
rect 941 -466 943 -452
rect 1008 -450 1010 -447
rect 1018 -450 1020 -447
rect 803 -494 805 -491
rect 745 -508 747 -499
rect 803 -520 805 -506
rect 842 -508 844 -481
rect 852 -508 854 -482
rect 870 -484 872 -473
rect 870 -508 872 -488
rect 880 -495 882 -473
rect 941 -475 943 -472
rect 980 -477 982 -468
rect 990 -478 992 -468
rect 941 -495 943 -492
rect 880 -508 882 -499
rect 707 -523 709 -520
rect 717 -523 719 -520
rect 735 -523 737 -520
rect 745 -523 747 -520
rect 842 -523 844 -520
rect 852 -523 854 -520
rect 870 -523 872 -520
rect 880 -523 882 -520
rect 941 -521 943 -507
rect 980 -509 982 -482
rect 990 -509 992 -483
rect 1008 -485 1010 -474
rect 1008 -509 1010 -489
rect 1018 -496 1020 -474
rect 1018 -509 1020 -500
rect 668 -529 670 -526
rect 803 -529 805 -526
rect 980 -524 982 -521
rect 990 -524 992 -521
rect 1008 -524 1010 -521
rect 1018 -524 1020 -521
rect 941 -530 943 -527
rect 567 -540 569 -537
rect 577 -540 579 -537
rect 595 -540 597 -537
rect 605 -540 607 -537
rect 528 -546 530 -543
rect 661 -568 663 -565
rect 697 -567 699 -564
rect 735 -567 737 -564
rect 455 -581 457 -578
rect 465 -581 467 -578
rect 497 -581 499 -578
rect 774 -568 776 -565
rect 455 -616 457 -593
rect 465 -616 467 -593
rect 497 -611 499 -593
rect 661 -595 663 -580
rect 697 -594 699 -579
rect 735 -594 737 -579
rect 823 -574 825 -571
rect 774 -595 776 -580
rect 890 -583 892 -580
rect 823 -604 825 -586
rect 929 -587 931 -584
rect 939 -587 941 -584
rect 890 -609 892 -595
rect 497 -621 499 -618
rect 553 -623 555 -615
rect 560 -623 562 -615
rect 607 -622 609 -615
rect 640 -622 642 -615
rect 671 -622 673 -615
rect 705 -621 707 -614
rect 726 -621 728 -614
rect 748 -621 750 -614
rect 776 -620 778 -613
rect 823 -614 825 -611
rect 957 -593 959 -590
rect 967 -593 969 -590
rect 890 -618 892 -615
rect 929 -620 931 -611
rect 455 -633 457 -629
rect 465 -633 467 -629
rect 455 -655 457 -652
rect 465 -655 467 -652
rect 497 -655 499 -652
rect 455 -690 457 -667
rect 465 -690 467 -667
rect 497 -685 499 -667
rect 497 -695 499 -692
rect 455 -707 457 -703
rect 465 -707 467 -703
rect 455 -724 457 -721
rect 465 -724 467 -721
rect 497 -724 499 -721
rect 455 -759 457 -736
rect 465 -759 467 -736
rect 497 -754 499 -736
rect 497 -764 499 -761
rect 455 -776 457 -772
rect 465 -776 467 -772
rect 455 -798 457 -795
rect 465 -798 467 -795
rect 497 -798 499 -795
rect 455 -833 457 -810
rect 465 -833 467 -810
rect 497 -828 499 -810
rect 497 -838 499 -835
rect 939 -621 941 -611
rect 890 -638 892 -635
rect 828 -650 830 -647
rect 828 -680 830 -662
rect 890 -664 892 -650
rect 929 -652 931 -625
rect 939 -652 941 -626
rect 957 -628 959 -617
rect 957 -652 959 -632
rect 967 -639 969 -617
rect 967 -652 969 -643
rect 929 -667 931 -664
rect 939 -667 941 -664
rect 957 -667 959 -664
rect 967 -667 969 -664
rect 890 -673 892 -670
rect 828 -690 830 -687
rect 901 -719 903 -716
rect 831 -726 833 -723
rect 940 -723 942 -720
rect 950 -723 952 -720
rect 831 -756 833 -738
rect 901 -745 903 -731
rect 968 -729 970 -726
rect 978 -729 980 -726
rect 901 -754 903 -751
rect 940 -756 942 -747
rect 950 -757 952 -747
rect 831 -766 833 -763
rect 901 -774 903 -771
rect 832 -798 834 -795
rect 901 -800 903 -786
rect 940 -788 942 -761
rect 950 -788 952 -762
rect 968 -764 970 -753
rect 968 -788 970 -768
rect 978 -775 980 -753
rect 978 -788 980 -779
rect 940 -803 942 -800
rect 950 -803 952 -800
rect 968 -803 970 -800
rect 978 -803 980 -800
rect 901 -809 903 -806
rect 832 -828 834 -810
rect 553 -839 555 -836
rect 560 -839 562 -836
rect 607 -839 609 -835
rect 640 -839 642 -835
rect 671 -839 673 -835
rect 705 -838 707 -834
rect 726 -838 728 -834
rect 748 -838 750 -834
rect 776 -837 778 -833
rect 832 -838 834 -835
rect 455 -850 457 -846
rect 465 -850 467 -846
rect 910 -853 912 -850
rect 949 -857 951 -854
rect 959 -857 961 -854
rect 910 -879 912 -865
rect 491 -884 493 -881
rect 977 -863 979 -860
rect 987 -863 989 -860
rect 910 -888 912 -885
rect 949 -890 951 -881
rect 959 -891 961 -881
rect 491 -914 493 -896
rect 910 -908 912 -905
rect 491 -924 493 -921
rect 910 -934 912 -920
rect 949 -922 951 -895
rect 959 -922 961 -896
rect 977 -898 979 -887
rect 977 -922 979 -902
rect 987 -909 989 -887
rect 987 -922 989 -913
rect 949 -937 951 -934
rect 959 -937 961 -934
rect 977 -937 979 -934
rect 987 -937 989 -934
rect 910 -943 912 -940
rect 340 -973 344 -971
rect 548 -973 555 -971
rect 915 -1002 917 -999
rect 954 -1006 956 -1003
rect 964 -1006 966 -1003
rect 915 -1028 917 -1014
rect 982 -1012 984 -1009
rect 992 -1012 994 -1009
rect 915 -1037 917 -1034
rect 954 -1039 956 -1030
rect 964 -1040 966 -1030
rect 915 -1057 917 -1054
rect 915 -1083 917 -1069
rect 954 -1071 956 -1044
rect 964 -1071 966 -1045
rect 982 -1047 984 -1036
rect 982 -1071 984 -1051
rect 992 -1058 994 -1036
rect 992 -1071 994 -1062
rect 954 -1086 956 -1083
rect 964 -1086 966 -1083
rect 982 -1086 984 -1083
rect 992 -1086 994 -1083
rect 915 -1092 917 -1089
<< polycontact >>
rect 524 -479 528 -475
rect 664 -462 668 -458
rect 799 -462 803 -458
rect 524 -534 528 -530
rect 593 -505 597 -501
rect 604 -516 608 -512
rect 664 -517 668 -513
rect 733 -488 737 -484
rect 937 -463 941 -459
rect 744 -499 748 -495
rect 799 -517 803 -513
rect 868 -488 872 -484
rect 879 -499 883 -495
rect 937 -518 941 -514
rect 1006 -489 1010 -485
rect 1017 -500 1021 -496
rect 451 -606 455 -602
rect 461 -613 465 -609
rect 493 -607 497 -603
rect 657 -595 661 -591
rect 693 -594 697 -590
rect 731 -594 735 -590
rect 770 -595 774 -591
rect 819 -600 823 -596
rect 886 -606 890 -602
rect 549 -619 553 -615
rect 562 -619 566 -615
rect 603 -619 607 -615
rect 636 -619 640 -615
rect 667 -619 671 -615
rect 701 -618 705 -614
rect 722 -618 726 -614
rect 744 -618 748 -614
rect 772 -617 776 -613
rect 451 -680 455 -676
rect 461 -687 465 -683
rect 493 -681 497 -677
rect 451 -749 455 -745
rect 461 -756 465 -752
rect 493 -750 497 -746
rect 451 -823 455 -819
rect 461 -830 465 -826
rect 493 -824 497 -820
rect 886 -661 890 -657
rect 824 -676 828 -672
rect 955 -632 959 -628
rect 966 -643 970 -639
rect 827 -752 831 -748
rect 897 -742 901 -738
rect 897 -797 901 -793
rect 966 -768 970 -764
rect 977 -779 981 -775
rect 828 -824 832 -820
rect 906 -876 910 -872
rect 487 -910 491 -906
rect 906 -931 910 -927
rect 975 -902 979 -898
rect 986 -913 990 -909
rect 551 -971 555 -967
rect 911 -1025 915 -1021
rect 911 -1080 915 -1076
rect 980 -1051 984 -1047
rect 991 -1062 995 -1058
<< metal1 >>
rect 662 -433 690 -430
rect 797 -433 825 -430
rect 663 -439 666 -433
rect 687 -434 690 -433
rect 687 -437 758 -434
rect 522 -450 550 -447
rect 523 -456 526 -450
rect 547 -451 550 -450
rect 547 -454 618 -451
rect 506 -480 509 -477
rect 514 -479 524 -476
rect 532 -476 535 -468
rect 562 -460 565 -454
rect 581 -460 584 -454
rect 532 -479 553 -476
rect 532 -482 535 -479
rect 523 -492 526 -488
rect 517 -494 541 -492
rect 517 -495 535 -494
rect 540 -495 541 -494
rect 550 -502 553 -479
rect 591 -460 611 -457
rect 591 -466 594 -460
rect 608 -466 611 -460
rect 646 -463 649 -460
rect 654 -462 664 -459
rect 672 -459 675 -451
rect 702 -443 705 -437
rect 721 -443 724 -437
rect 798 -439 801 -433
rect 822 -434 825 -433
rect 935 -434 963 -431
rect 822 -437 893 -434
rect 672 -462 693 -459
rect 672 -465 675 -462
rect 572 -487 575 -484
rect 572 -490 590 -487
rect 663 -475 666 -471
rect 657 -477 681 -475
rect 657 -478 675 -477
rect 680 -478 681 -477
rect 690 -485 693 -462
rect 731 -443 751 -440
rect 731 -449 734 -443
rect 748 -449 751 -443
rect 712 -470 715 -467
rect 712 -473 730 -470
rect 781 -463 784 -460
rect 789 -462 799 -459
rect 807 -459 810 -451
rect 837 -443 840 -437
rect 856 -443 859 -437
rect 936 -440 939 -434
rect 960 -435 963 -434
rect 960 -438 1031 -435
rect 807 -462 828 -459
rect 807 -465 810 -462
rect 740 -480 743 -473
rect 798 -475 801 -471
rect 792 -477 816 -475
rect 792 -478 810 -477
rect 740 -483 757 -480
rect 662 -486 681 -485
rect 657 -488 681 -486
rect 690 -488 733 -485
rect 600 -497 603 -490
rect 663 -494 666 -488
rect 754 -494 757 -483
rect 815 -478 816 -477
rect 825 -485 828 -462
rect 866 -443 886 -440
rect 866 -449 869 -443
rect 883 -449 886 -443
rect 847 -470 850 -467
rect 847 -473 865 -470
rect 919 -464 922 -461
rect 927 -463 937 -460
rect 945 -460 948 -452
rect 975 -444 978 -438
rect 994 -444 997 -438
rect 945 -463 966 -460
rect 945 -466 948 -463
rect 875 -480 878 -473
rect 936 -476 939 -472
rect 930 -478 954 -476
rect 930 -479 948 -478
rect 875 -483 892 -480
rect 797 -486 816 -485
rect 792 -488 816 -486
rect 825 -488 868 -485
rect 798 -494 801 -488
rect 889 -494 892 -483
rect 953 -479 954 -478
rect 963 -486 966 -463
rect 1004 -444 1024 -441
rect 1004 -450 1007 -444
rect 1021 -450 1024 -444
rect 985 -471 988 -468
rect 985 -474 1003 -471
rect 1013 -481 1016 -474
rect 1013 -484 1030 -481
rect 935 -487 954 -486
rect 930 -489 954 -487
rect 963 -489 1006 -486
rect 600 -500 617 -497
rect 522 -503 541 -502
rect 517 -505 541 -503
rect 550 -505 593 -502
rect 523 -511 526 -505
rect 614 -511 617 -500
rect 719 -499 744 -496
rect 754 -498 766 -494
rect 719 -501 722 -499
rect 579 -516 604 -513
rect 614 -515 627 -511
rect 579 -518 582 -516
rect 506 -534 509 -531
rect 514 -534 524 -531
rect 532 -531 535 -523
rect 544 -521 582 -518
rect 614 -519 617 -515
rect 544 -531 547 -521
rect 585 -522 617 -519
rect 585 -525 588 -522
rect 532 -534 547 -531
rect 532 -537 535 -534
rect 584 -528 590 -525
rect 523 -547 526 -543
rect 544 -544 549 -541
rect 562 -541 565 -537
rect 609 -541 612 -537
rect 554 -544 618 -541
rect 544 -547 547 -544
rect 517 -550 547 -547
rect 623 -548 627 -515
rect 646 -517 649 -514
rect 654 -517 664 -514
rect 672 -514 675 -506
rect 684 -504 722 -501
rect 754 -502 757 -498
rect 684 -514 687 -504
rect 725 -505 757 -502
rect 725 -508 728 -505
rect 672 -517 687 -514
rect 672 -520 675 -517
rect 724 -511 730 -508
rect 663 -530 666 -526
rect 684 -527 689 -524
rect 702 -524 705 -520
rect 749 -524 752 -520
rect 694 -527 758 -524
rect 684 -530 687 -527
rect 657 -533 687 -530
rect 762 -534 766 -498
rect 854 -499 879 -496
rect 889 -498 900 -494
rect 854 -501 857 -499
rect 781 -517 784 -514
rect 789 -517 799 -514
rect 807 -514 810 -506
rect 819 -504 857 -501
rect 889 -502 892 -498
rect 819 -514 822 -504
rect 860 -505 892 -502
rect 860 -508 863 -505
rect 807 -517 822 -514
rect 807 -520 810 -517
rect 859 -511 865 -508
rect 798 -530 801 -526
rect 819 -527 824 -524
rect 837 -524 840 -520
rect 884 -524 887 -520
rect 829 -527 893 -524
rect 819 -530 822 -527
rect 792 -533 822 -530
rect 702 -537 766 -534
rect 568 -552 627 -548
rect 633 -538 766 -537
rect 896 -538 900 -498
rect 936 -495 939 -489
rect 1027 -495 1030 -484
rect 992 -500 1017 -497
rect 1027 -499 1042 -495
rect 992 -502 995 -500
rect 919 -518 922 -515
rect 927 -518 937 -515
rect 945 -515 948 -507
rect 957 -505 995 -502
rect 1027 -503 1030 -499
rect 957 -515 960 -505
rect 998 -506 1030 -503
rect 998 -509 1001 -506
rect 945 -518 960 -515
rect 945 -521 948 -518
rect 997 -512 1003 -509
rect 936 -531 939 -527
rect 957 -528 962 -525
rect 975 -525 978 -521
rect 1022 -525 1025 -521
rect 967 -528 1031 -525
rect 957 -531 960 -528
rect 930 -534 960 -531
rect 1038 -535 1042 -499
rect 633 -541 706 -538
rect 442 -575 513 -572
rect 450 -581 454 -575
rect 468 -581 472 -575
rect 492 -581 495 -575
rect 459 -596 462 -593
rect 459 -599 472 -596
rect 436 -602 442 -601
rect 436 -606 451 -602
rect 469 -603 472 -599
rect 501 -603 504 -593
rect 469 -607 493 -603
rect 501 -606 513 -603
rect 442 -613 461 -609
rect 469 -616 472 -607
rect 501 -611 504 -606
rect 568 -608 572 -552
rect 633 -555 637 -541
rect 773 -542 900 -538
rect 710 -546 777 -542
rect 643 -550 714 -546
rect 643 -552 647 -550
rect 587 -559 637 -555
rect 640 -556 647 -552
rect 568 -612 575 -608
rect 571 -615 575 -612
rect 450 -635 453 -629
rect 492 -635 495 -618
rect 546 -619 549 -615
rect 566 -619 575 -615
rect 587 -615 591 -559
rect 640 -581 644 -556
rect 649 -562 677 -559
rect 685 -561 713 -558
rect 723 -561 751 -558
rect 656 -568 659 -562
rect 692 -567 695 -561
rect 730 -567 733 -561
rect 762 -562 790 -559
rect 625 -585 644 -581
rect 625 -615 629 -585
rect 649 -595 657 -591
rect 665 -608 668 -580
rect 685 -594 693 -590
rect 701 -601 704 -579
rect 723 -594 731 -590
rect 701 -604 724 -601
rect 721 -608 724 -604
rect 739 -606 742 -579
rect 769 -568 772 -562
rect 811 -568 843 -565
rect 762 -595 770 -591
rect 778 -594 781 -580
rect 818 -574 821 -568
rect 884 -577 912 -574
rect 665 -611 712 -608
rect 721 -611 733 -608
rect 739 -610 755 -606
rect 778 -607 782 -594
rect 827 -596 830 -586
rect 885 -583 888 -577
rect 909 -578 912 -577
rect 909 -581 980 -578
rect 807 -600 819 -596
rect 827 -599 839 -596
rect 827 -604 830 -599
rect 709 -614 712 -611
rect 587 -619 603 -615
rect 625 -619 636 -615
rect 664 -619 667 -615
rect 674 -622 678 -615
rect 698 -618 701 -614
rect 708 -621 712 -614
rect 719 -618 722 -614
rect 729 -621 733 -611
rect 741 -618 744 -614
rect 751 -621 755 -610
rect 769 -617 772 -613
rect 779 -620 783 -607
rect 442 -638 495 -635
rect 442 -649 513 -646
rect 450 -655 454 -649
rect 468 -655 472 -649
rect 492 -655 495 -649
rect 459 -670 462 -667
rect 459 -673 472 -670
rect 436 -676 442 -675
rect 436 -680 451 -676
rect 469 -677 472 -673
rect 501 -677 504 -667
rect 469 -681 493 -677
rect 501 -680 513 -677
rect 442 -687 461 -683
rect 469 -690 472 -681
rect 501 -685 504 -680
rect 450 -709 453 -703
rect 492 -709 495 -692
rect 442 -712 495 -709
rect 442 -718 513 -715
rect 450 -724 454 -718
rect 468 -724 472 -718
rect 492 -724 495 -718
rect 459 -739 462 -736
rect 459 -742 472 -739
rect 436 -749 451 -745
rect 469 -746 472 -742
rect 501 -746 504 -736
rect 469 -750 493 -746
rect 501 -749 513 -746
rect 442 -756 461 -752
rect 469 -759 472 -750
rect 501 -754 504 -749
rect 450 -778 453 -772
rect 492 -778 495 -761
rect 442 -781 495 -778
rect 442 -792 513 -789
rect 450 -798 454 -792
rect 468 -798 472 -792
rect 492 -798 495 -792
rect 459 -813 462 -810
rect 459 -816 472 -813
rect 436 -823 451 -819
rect 469 -820 472 -816
rect 501 -820 504 -810
rect 469 -824 493 -820
rect 501 -823 513 -820
rect 442 -830 461 -826
rect 469 -833 472 -824
rect 501 -828 504 -823
rect 450 -852 453 -846
rect 492 -852 495 -835
rect 548 -845 552 -836
rect 563 -837 568 -836
rect 602 -837 606 -835
rect 563 -842 606 -837
rect 610 -837 614 -835
rect 635 -837 639 -835
rect 610 -842 639 -837
rect 643 -837 647 -835
rect 868 -607 871 -604
rect 876 -606 886 -603
rect 894 -603 897 -595
rect 924 -587 927 -581
rect 943 -587 946 -581
rect 894 -606 915 -603
rect 894 -609 897 -606
rect 818 -628 821 -611
rect 885 -619 888 -615
rect 879 -621 903 -619
rect 879 -622 897 -621
rect 807 -631 821 -628
rect 902 -622 903 -621
rect 912 -629 915 -606
rect 953 -587 973 -584
rect 953 -593 956 -587
rect 970 -593 973 -587
rect 934 -614 937 -611
rect 934 -617 952 -614
rect 962 -624 965 -617
rect 962 -627 979 -624
rect 884 -630 903 -629
rect 879 -632 903 -630
rect 912 -632 955 -629
rect 885 -638 888 -632
rect 976 -638 979 -627
rect 1003 -638 1019 -635
rect 812 -644 844 -641
rect 823 -650 826 -644
rect 976 -639 1019 -638
rect 941 -643 966 -640
rect 976 -642 1007 -639
rect 941 -645 944 -643
rect 868 -661 871 -658
rect 876 -661 886 -658
rect 894 -658 897 -650
rect 906 -648 944 -645
rect 976 -646 979 -642
rect 906 -658 909 -648
rect 947 -649 979 -646
rect 947 -652 950 -649
rect 894 -661 909 -658
rect 832 -672 835 -662
rect 894 -664 897 -661
rect 946 -655 952 -652
rect 812 -676 824 -672
rect 832 -675 844 -672
rect 885 -674 888 -670
rect 906 -671 911 -668
rect 924 -668 927 -664
rect 971 -668 974 -664
rect 916 -671 980 -668
rect 906 -674 909 -671
rect 832 -680 835 -675
rect 879 -677 909 -674
rect 823 -704 826 -687
rect 812 -707 826 -704
rect 895 -713 923 -710
rect 815 -720 847 -717
rect 896 -719 899 -713
rect 920 -714 923 -713
rect 920 -717 991 -714
rect 826 -726 829 -720
rect 835 -748 838 -738
rect 879 -743 882 -740
rect 887 -742 897 -739
rect 905 -739 908 -731
rect 935 -723 938 -717
rect 954 -723 957 -717
rect 905 -742 926 -739
rect 905 -745 908 -742
rect 815 -752 827 -748
rect 835 -751 847 -748
rect 835 -756 838 -751
rect 896 -755 899 -751
rect 890 -757 914 -755
rect 890 -758 908 -757
rect 826 -780 829 -763
rect 913 -758 914 -757
rect 923 -765 926 -742
rect 964 -723 984 -720
rect 964 -729 967 -723
rect 981 -729 984 -723
rect 945 -750 948 -747
rect 945 -753 963 -750
rect 973 -760 976 -753
rect 973 -763 990 -760
rect 895 -766 914 -765
rect 890 -768 914 -766
rect 923 -768 966 -765
rect 815 -783 829 -780
rect 896 -774 899 -768
rect 987 -774 990 -763
rect 952 -779 977 -776
rect 987 -778 1019 -774
rect 952 -781 955 -779
rect 816 -792 848 -789
rect 827 -798 830 -792
rect 879 -797 882 -794
rect 887 -797 897 -794
rect 905 -794 908 -786
rect 917 -784 955 -781
rect 987 -782 990 -778
rect 917 -794 920 -784
rect 958 -785 990 -782
rect 958 -788 961 -785
rect 905 -797 920 -794
rect 905 -800 908 -797
rect 957 -791 963 -788
rect 896 -810 899 -806
rect 917 -807 922 -804
rect 935 -804 938 -800
rect 982 -804 985 -800
rect 927 -807 991 -804
rect 917 -810 920 -807
rect 836 -820 839 -810
rect 890 -813 920 -810
rect 816 -824 828 -820
rect 836 -823 848 -820
rect 836 -828 839 -823
rect 666 -837 670 -835
rect 643 -842 670 -837
rect 700 -839 704 -834
rect 721 -839 725 -834
rect 743 -839 747 -834
rect 771 -839 775 -833
rect 700 -842 775 -839
rect 543 -849 561 -845
rect 827 -852 830 -835
rect 904 -847 932 -844
rect 442 -855 495 -852
rect 816 -855 830 -852
rect 905 -853 908 -847
rect 929 -848 932 -847
rect 929 -851 1000 -848
rect 476 -878 507 -875
rect 888 -877 891 -874
rect 896 -876 906 -873
rect 914 -873 917 -865
rect 944 -857 947 -851
rect 963 -857 966 -851
rect 914 -876 935 -873
rect 486 -884 489 -878
rect 914 -879 917 -876
rect 905 -889 908 -885
rect 899 -891 923 -889
rect 899 -892 917 -891
rect 495 -906 498 -896
rect 922 -892 923 -891
rect 932 -899 935 -876
rect 973 -857 993 -854
rect 973 -863 976 -857
rect 990 -863 993 -857
rect 954 -884 957 -881
rect 954 -887 972 -884
rect 982 -894 985 -887
rect 982 -897 999 -894
rect 904 -900 923 -899
rect 899 -902 923 -900
rect 932 -902 975 -899
rect 476 -910 487 -906
rect 495 -909 507 -906
rect 905 -908 908 -902
rect 996 -908 999 -897
rect 495 -914 498 -909
rect 961 -913 986 -910
rect 996 -912 1019 -908
rect 961 -915 964 -913
rect 486 -938 489 -921
rect 888 -931 891 -928
rect 896 -931 906 -928
rect 914 -928 917 -920
rect 926 -918 964 -915
rect 996 -916 999 -912
rect 926 -928 929 -918
rect 967 -919 999 -916
rect 967 -922 970 -919
rect 914 -931 929 -928
rect 914 -934 917 -931
rect 476 -941 489 -938
rect 966 -925 972 -922
rect 905 -944 908 -940
rect 926 -941 931 -938
rect 944 -938 947 -934
rect 991 -938 994 -934
rect 936 -941 1000 -938
rect 926 -944 929 -941
rect 899 -947 929 -944
rect 337 -966 342 -958
rect 337 -970 344 -966
rect 551 -967 555 -958
rect 337 -978 344 -974
rect 337 -985 342 -978
rect 909 -996 937 -993
rect 910 -1002 913 -996
rect 934 -997 937 -996
rect 934 -1000 1005 -997
rect 893 -1026 896 -1023
rect 901 -1025 911 -1022
rect 919 -1022 922 -1014
rect 949 -1006 952 -1000
rect 968 -1006 971 -1000
rect 919 -1025 940 -1022
rect 919 -1028 922 -1025
rect 910 -1038 913 -1034
rect 904 -1040 928 -1038
rect 904 -1041 922 -1040
rect 927 -1041 928 -1040
rect 937 -1048 940 -1025
rect 978 -1006 998 -1003
rect 978 -1012 981 -1006
rect 995 -1012 998 -1006
rect 959 -1033 962 -1030
rect 959 -1036 977 -1033
rect 987 -1043 990 -1036
rect 987 -1046 1004 -1043
rect 909 -1049 928 -1048
rect 904 -1051 928 -1049
rect 937 -1051 980 -1048
rect 910 -1057 913 -1051
rect 1001 -1057 1004 -1046
rect 966 -1062 991 -1059
rect 1001 -1061 1019 -1057
rect 966 -1064 969 -1062
rect 893 -1080 896 -1077
rect 901 -1080 911 -1077
rect 919 -1077 922 -1069
rect 931 -1067 969 -1064
rect 1001 -1065 1004 -1061
rect 931 -1077 934 -1067
rect 972 -1068 1004 -1065
rect 972 -1071 975 -1068
rect 919 -1080 934 -1077
rect 919 -1083 922 -1080
rect 971 -1074 977 -1071
rect 910 -1093 913 -1089
rect 931 -1090 936 -1087
rect 949 -1087 952 -1083
rect 996 -1087 999 -1083
rect 941 -1090 1005 -1087
rect 931 -1093 934 -1090
rect 904 -1096 934 -1093
<< m2contact >>
rect 509 -481 514 -476
rect 649 -464 654 -459
rect 784 -464 789 -459
rect 922 -465 927 -460
rect 509 -535 514 -530
rect 649 -518 654 -513
rect 784 -518 789 -513
rect 922 -519 927 -514
rect 668 -599 673 -594
rect 724 -608 729 -603
rect 802 -600 807 -595
rect 755 -617 760 -612
rect 871 -608 876 -603
rect 871 -662 876 -657
rect 807 -676 812 -671
rect 810 -752 815 -747
rect 882 -744 887 -739
rect 882 -798 887 -793
rect 891 -878 896 -873
rect 891 -932 896 -927
rect 896 -1027 901 -1022
rect 896 -1081 901 -1076
<< pm12contact >>
rect 705 -481 710 -476
rect 714 -482 719 -477
rect 565 -498 570 -493
rect 574 -499 579 -494
rect 840 -481 845 -476
rect 849 -482 854 -477
rect 978 -482 983 -477
rect 987 -483 992 -478
rect 927 -625 932 -620
rect 936 -626 941 -621
rect 938 -761 943 -756
rect 947 -762 952 -757
rect 947 -895 952 -890
rect 956 -896 961 -891
rect 952 -1044 957 -1039
rect 961 -1045 966 -1040
<< metal2 >>
rect 650 -470 653 -464
rect 785 -470 788 -464
rect 650 -473 687 -470
rect 785 -473 822 -470
rect 684 -476 687 -473
rect 819 -476 822 -473
rect 923 -471 926 -465
rect 923 -474 960 -471
rect 510 -487 513 -481
rect 684 -479 705 -476
rect 510 -490 547 -487
rect 544 -493 547 -490
rect 714 -492 717 -482
rect 819 -479 840 -476
rect 957 -477 960 -474
rect 849 -492 852 -482
rect 957 -480 978 -477
rect 544 -496 565 -493
rect 651 -495 717 -492
rect 786 -495 852 -492
rect 987 -493 990 -483
rect 574 -509 577 -499
rect 511 -512 577 -509
rect 511 -530 514 -512
rect 651 -513 654 -495
rect 786 -513 789 -495
rect 924 -496 990 -493
rect 924 -514 927 -496
rect 673 -599 802 -595
rect 729 -608 806 -604
rect 755 -620 760 -617
rect 756 -752 759 -620
rect 802 -669 806 -608
rect 872 -614 875 -608
rect 872 -617 909 -614
rect 906 -620 909 -617
rect 906 -623 927 -620
rect 936 -636 939 -626
rect 873 -639 939 -636
rect 873 -657 876 -639
rect 802 -672 807 -669
rect 804 -676 807 -672
rect 806 -752 810 -747
rect 883 -750 886 -744
rect 756 -755 810 -752
rect 883 -753 920 -750
rect 917 -756 920 -753
rect 917 -759 938 -756
rect 947 -772 950 -762
rect 884 -775 950 -772
rect 884 -793 887 -775
rect 916 -790 919 -787
rect 892 -884 895 -878
rect 892 -887 929 -884
rect 926 -890 929 -887
rect 926 -893 947 -890
rect 956 -906 959 -896
rect 893 -909 959 -906
rect 893 -927 896 -909
rect 897 -1033 900 -1027
rect 897 -1036 934 -1033
rect 931 -1039 934 -1036
rect 931 -1042 952 -1039
rect 961 -1055 964 -1045
rect 898 -1058 964 -1055
rect 898 -1076 901 -1058
<< m3contact >>
rect 1038 -540 1043 -535
rect 513 -608 518 -603
rect 437 -613 442 -608
rect 659 -619 664 -614
rect 693 -618 698 -613
rect 714 -618 719 -613
rect 736 -618 741 -613
rect 764 -617 769 -612
rect 783 -620 788 -614
rect 513 -682 518 -677
rect 437 -687 442 -682
rect 513 -751 518 -746
rect 437 -756 442 -751
rect 513 -825 518 -820
rect 811 -824 816 -819
rect 437 -830 442 -825
<< m123contact >>
rect 657 -433 662 -428
rect 792 -433 797 -428
rect 930 -434 935 -429
rect 517 -450 522 -445
rect 657 -486 662 -481
rect 675 -482 680 -477
rect 792 -486 797 -481
rect 810 -482 815 -477
rect 930 -487 935 -482
rect 948 -483 953 -478
rect 517 -503 522 -498
rect 535 -499 540 -494
rect 689 -527 694 -522
rect 824 -527 829 -522
rect 962 -528 967 -523
rect 549 -544 554 -539
rect 879 -577 884 -572
rect 879 -630 884 -625
rect 897 -626 902 -621
rect 911 -671 916 -666
rect 890 -713 895 -708
rect 890 -766 895 -761
rect 908 -762 913 -757
rect 922 -807 927 -802
rect 899 -847 904 -842
rect 899 -900 904 -895
rect 917 -896 922 -891
rect 931 -941 936 -936
rect 904 -996 909 -991
rect 904 -1049 909 -1044
rect 922 -1045 927 -1040
rect 936 -1090 941 -1085
<< metal3 >>
rect 517 -498 520 -450
rect 657 -481 660 -433
rect 680 -482 692 -479
rect 540 -499 552 -496
rect 549 -539 552 -499
rect 689 -522 692 -482
rect 792 -481 795 -433
rect 815 -482 827 -479
rect 824 -522 827 -482
rect 930 -482 933 -434
rect 953 -483 965 -480
rect 962 -523 965 -483
rect 975 -540 1038 -535
rect 975 -544 980 -540
rect 911 -549 980 -544
rect 911 -553 916 -549
rect 631 -558 916 -553
rect 631 -596 636 -558
rect 631 -601 648 -596
rect 518 -608 535 -603
rect 436 -613 437 -608
rect 530 -639 535 -608
rect 643 -604 648 -601
rect 643 -609 657 -604
rect 652 -614 657 -609
rect 652 -619 659 -614
rect 687 -618 693 -613
rect 687 -639 692 -618
rect 714 -623 718 -618
rect 530 -644 692 -639
rect 713 -677 718 -623
rect 518 -682 718 -677
rect 436 -687 437 -682
rect 736 -746 741 -618
rect 518 -751 741 -746
rect 760 -617 764 -612
rect 436 -756 437 -751
rect 760 -820 765 -617
rect 518 -825 765 -820
rect 788 -819 793 -614
rect 879 -625 882 -577
rect 902 -626 914 -623
rect 911 -666 914 -626
rect 890 -761 893 -713
rect 913 -762 925 -759
rect 922 -802 925 -762
rect 788 -824 811 -819
rect 788 -825 793 -824
rect 436 -830 437 -825
rect 899 -895 902 -847
rect 922 -896 934 -893
rect 931 -936 934 -896
rect 904 -1044 907 -996
rect 927 -1045 939 -1042
rect 936 -1085 939 -1045
<< labels >>
rlabel metal1 535 -550 539 -547 1 gnd
rlabel metal1 585 -544 588 -542 1 gnd
rlabel metal1 533 -494 534 -492 1 gnd
rlabel metal1 529 -450 532 -448 5 vdd
rlabel metal1 530 -504 533 -502 1 vdd
rlabel metal1 614 -515 618 -511 7 p0
rlabel metal1 506 -480 507 -477 1 a0
rlabel metal1 506 -534 507 -531 1 b0
rlabel metal1 508 -605 509 -604 7 g0
rlabel metal1 445 -611 446 -610 3 b0
rlabel metal1 443 -604 444 -603 3 a0
rlabel metal1 468 -637 468 -637 1 gnd!
rlabel metal1 468 -573 468 -573 5 vdd!
rlabel metal1 508 -679 509 -678 7 g1
rlabel metal1 468 -780 468 -780 1 gnd!
rlabel metal1 468 -716 468 -716 5 vdd!
rlabel metal1 468 -854 468 -854 1 gnd!
rlabel metal1 468 -790 468 -790 5 vdd!
rlabel metal1 443 -747 444 -746 3 a2
rlabel metal1 445 -754 446 -753 3 b2
rlabel metal1 444 -821 445 -820 3 a3
rlabel metal1 445 -828 446 -827 3 b3
rlabel metal1 508 -822 509 -821 7 g3
rlabel metal1 445 -685 446 -684 3 b1
rlabel metal1 444 -678 445 -677 3 a1
rlabel metal1 468 -647 468 -647 5 vdd!
rlabel metal1 468 -711 468 -711 1 gnd!
rlabel metal1 547 -618 548 -617 1 cin
rlabel metal1 568 -618 569 -616 1 p0
rlabel metal1 601 -618 602 -617 1 p1
rlabel metal1 634 -618 635 -617 1 p2
rlabel metal1 665 -618 666 -617 1 p3
rlabel metal1 675 -619 677 -617 1 c3b
rlabel metal1 699 -617 700 -616 1 g0
rlabel metal1 709 -618 711 -616 1 c0b
rlabel metal1 720 -617 721 -616 1 g1
rlabel metal1 730 -618 732 -616 1 c1b
rlabel metal1 897 -677 901 -674 1 gnd
rlabel metal1 947 -671 950 -669 1 gnd
rlabel metal1 895 -621 896 -619 1 gnd
rlabel metal1 891 -577 894 -575 5 vdd
rlabel metal1 892 -631 895 -629 1 vdd
rlabel metal1 908 -813 912 -810 1 gnd
rlabel metal1 958 -807 961 -805 1 gnd
rlabel metal1 906 -757 907 -755 1 gnd
rlabel metal1 902 -713 905 -711 5 vdd
rlabel metal1 903 -767 906 -765 1 vdd
rlabel metal1 917 -947 921 -944 1 gnd
rlabel metal1 967 -941 970 -939 1 gnd
rlabel metal1 915 -891 916 -889 1 gnd
rlabel metal1 911 -847 914 -845 5 vdd
rlabel metal1 912 -901 915 -899 1 vdd
rlabel metal1 922 -1096 926 -1093 1 gnd
rlabel metal1 972 -1090 975 -1088 1 gnd
rlabel metal1 920 -1040 921 -1038 1 gnd
rlabel metal1 916 -996 919 -994 5 vdd
rlabel metal1 917 -1050 920 -1048 1 vdd
rlabel metal1 868 -607 869 -604 1 p0
rlabel metal1 868 -661 869 -658 1 cin
rlabel metal1 976 -642 980 -638 1 s0
rlabel metal1 879 -743 880 -740 1 p1
rlabel metal1 879 -797 880 -794 1 c0
rlabel metal1 987 -778 991 -774 1 s1
rlabel metal1 888 -877 889 -874 1 p2
rlabel metal1 888 -931 889 -928 1 c1
rlabel metal1 996 -912 1000 -908 1 s2
rlabel metal1 893 -1026 894 -1023 1 p3
rlabel metal1 893 -1080 894 -1077 1 c2
rlabel metal1 1001 -1061 1005 -1057 1 s3
rlabel metal1 508 -748 509 -747 7 g2
rlabel metal1 662 -561 669 -560 1 vdd
rlabel metal1 666 -593 667 -592 1 c0b
rlabel metal1 702 -592 703 -591 1 c1b
rlabel metal1 698 -560 705 -559 1 vdd
rlabel metal1 736 -560 743 -559 1 vdd
rlabel metal1 740 -592 741 -591 1 c2b
rlabel metal1 675 -533 679 -530 1 gnd
rlabel metal1 725 -527 728 -525 1 gnd
rlabel metal1 673 -477 674 -475 1 gnd
rlabel metal1 669 -433 672 -431 5 vdd
rlabel metal1 670 -487 673 -485 1 vdd
rlabel metal1 810 -533 814 -530 1 gnd
rlabel metal1 860 -527 863 -525 1 gnd
rlabel metal1 808 -477 809 -475 1 gnd
rlabel metal1 804 -433 807 -431 5 vdd
rlabel metal1 805 -487 808 -485 1 vdd
rlabel metal1 948 -534 952 -531 1 gnd
rlabel metal1 998 -528 1001 -526 1 gnd
rlabel metal1 946 -478 947 -476 1 gnd
rlabel metal1 942 -434 945 -432 5 vdd
rlabel metal1 943 -488 946 -486 1 vdd
rlabel metal1 646 -517 647 -514 1 b1
rlabel metal1 646 -463 647 -460 1 a1
rlabel metal1 781 -463 782 -460 1 a2
rlabel metal1 781 -517 782 -514 1 b2
rlabel metal1 919 -464 920 -461 1 a3
rlabel metal1 919 -518 920 -515 1 b3
rlabel metal1 1027 -499 1031 -495 7 p3
rlabel metal1 754 -498 758 -494 1 p1
rlabel metal1 889 -498 893 -494 1 p2
rlabel metal1 770 -616 771 -615 1 g3
rlabel metal1 780 -617 782 -615 1 c3b
rlabel metal1 742 -617 743 -616 1 g2
rlabel metal1 752 -618 754 -616 1 c2b
rlabel metal1 816 -675 819 -673 1 c1b
rlabel metal1 839 -674 840 -673 1 c1
rlabel metal1 818 -706 820 -705 1 gnd
rlabel metal1 826 -643 828 -642 1 vdd
rlabel metal1 810 -599 811 -597 1 c0b
rlabel metal1 834 -598 837 -596 1 c0
rlabel metal1 811 -630 813 -629 1 gnd
rlabel metal1 820 -567 822 -566 1 vdd
rlabel metal1 775 -561 782 -560 1 vdd
rlabel metal1 779 -593 780 -592 1 c3b
rlabel metal1 820 -751 823 -749 1 c2b
rlabel metal1 821 -823 824 -821 1 c3b
rlabel metal1 842 -750 843 -749 1 c2
rlabel metal1 843 -822 844 -821 1 c3
rlabel metal1 821 -854 823 -853 1 gnd
rlabel metal1 828 -791 830 -790 1 vdd
rlabel metal1 821 -781 823 -780 1 gnd
rlabel metal1 827 -719 829 -718 1 vdd
rlabel metal1 651 -594 655 -592 1 clkb
rlabel metal1 687 -593 691 -591 1 clkb
rlabel metal1 724 -593 729 -591 1 clkb
rlabel metal1 763 -595 768 -592 1 clkb
rlabel metal1 552 -966 554 -964 1 clkb
rlabel metal1 338 -966 341 -960 1 k
rlabel metal1 338 -982 340 -977 1 gnd
rlabel metal1 480 -940 481 -939 1 gnd
rlabel metal1 490 -877 491 -876 1 vdd
rlabel metal1 502 -908 503 -907 1 clkb
rlabel metal1 480 -908 481 -907 1 clk
rlabel metal1 654 -842 661 -837 1 c2b
rlabel metal1 619 -842 626 -837 1 c1b
rlabel metal1 580 -842 587 -837 1 c0b
rlabel metal1 722 -842 727 -840 1 k
rlabel metal1 551 -848 559 -846 1 k
<< end >>
