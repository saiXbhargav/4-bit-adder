magic
tech scmos
timestamp 1732080275
<< nwell >>
rect 2638 684 2662 708
rect 2677 698 2711 704
rect 2778 701 2802 725
rect 2817 715 2851 721
rect 2186 641 2218 678
rect 2224 641 2250 678
rect 2268 641 2294 678
rect 2313 641 2339 678
rect 2381 644 2413 681
rect 2419 644 2445 681
rect 2463 644 2489 681
rect 2508 644 2534 681
rect 2677 668 2739 698
rect 2817 685 2879 715
rect 2913 701 2937 725
rect 2952 715 2986 721
rect 2952 685 3014 715
rect 3051 700 3075 724
rect 3090 714 3124 720
rect 2845 679 2879 685
rect 2980 679 3014 685
rect 3090 684 3152 714
rect 3118 678 3152 684
rect 2705 662 2739 668
rect 2638 629 2662 653
rect 2778 646 2802 670
rect 2913 646 2937 670
rect 3051 645 3075 669
rect 2183 540 2215 577
rect 2221 540 2247 577
rect 2265 540 2291 577
rect 2310 540 2336 577
rect 2383 546 2415 583
rect 2421 546 2447 583
rect 2465 546 2491 583
rect 2510 546 2536 583
rect 2563 557 2600 583
rect 2606 557 2634 583
rect 2770 570 2798 596
rect 2806 571 2834 597
rect 2844 571 2872 597
rect 2883 570 2911 596
rect 2932 564 2960 590
rect 3000 557 3024 581
rect 3039 571 3073 577
rect 3039 541 3101 571
rect 3067 535 3101 541
rect 2182 443 2214 480
rect 2220 443 2246 480
rect 2264 443 2290 480
rect 2309 443 2335 480
rect 2382 449 2414 486
rect 2420 449 2446 486
rect 2464 449 2490 486
rect 2509 449 2535 486
rect 2563 483 2600 509
rect 2606 483 2634 509
rect 2937 488 2965 514
rect 3000 502 3024 526
rect 3158 524 3190 561
rect 3196 524 3222 561
rect 3240 524 3266 561
rect 3285 524 3311 561
rect 2563 414 2600 440
rect 2606 414 2634 440
rect 2940 412 2968 438
rect 3011 421 3035 445
rect 3050 435 3084 441
rect 3050 405 3112 435
rect 3078 399 3112 405
rect 2183 347 2215 384
rect 2221 347 2247 384
rect 2265 347 2291 384
rect 2310 347 2336 384
rect 2383 353 2415 390
rect 2421 353 2447 390
rect 2465 353 2491 390
rect 2510 353 2536 390
rect 3011 366 3035 390
rect 3171 382 3203 419
rect 3209 382 3235 419
rect 3253 382 3279 419
rect 3298 382 3324 419
rect 2563 340 2600 366
rect 2606 340 2634 366
rect 2929 340 2957 366
rect 2385 252 2417 289
rect 2423 252 2449 289
rect 2467 252 2493 289
rect 2512 252 2538 289
rect 3020 287 3044 311
rect 3059 301 3093 307
rect 3059 271 3121 301
rect 3087 265 3121 271
rect 3181 259 3213 296
rect 3219 259 3245 296
rect 3263 259 3289 296
rect 3308 259 3334 296
rect 2731 198 2757 235
rect 2776 198 2802 235
rect 2820 198 2846 235
rect 2852 198 2884 235
rect 3020 232 3044 256
rect 3025 138 3049 162
rect 3064 152 3098 158
rect 3064 122 3126 152
rect 3092 116 3126 122
rect 3186 112 3218 149
rect 3224 112 3250 149
rect 3268 112 3294 149
rect 3313 112 3339 149
rect 3025 83 3049 107
<< ntransistor >>
rect 2649 670 2651 676
rect 2789 687 2791 693
rect 2924 687 2926 693
rect 2193 615 2195 625
rect 2229 615 2231 625
rect 2237 615 2239 625
rect 2273 615 2275 625
rect 2281 615 2283 625
rect 2324 615 2326 625
rect 2388 618 2390 628
rect 2424 618 2426 628
rect 2432 618 2434 628
rect 2468 618 2470 628
rect 2476 618 2478 628
rect 2519 618 2521 628
rect 3062 686 3064 692
rect 2828 638 2830 650
rect 2838 638 2840 650
rect 2856 638 2858 650
rect 2866 638 2868 650
rect 2963 638 2965 650
rect 2973 638 2975 650
rect 2991 638 2993 650
rect 3001 638 3003 650
rect 2688 621 2690 633
rect 2698 621 2700 633
rect 2716 621 2718 633
rect 2726 621 2728 633
rect 2789 632 2791 638
rect 2924 632 2926 638
rect 3101 637 3103 649
rect 3111 637 3113 649
rect 3129 637 3131 649
rect 3139 637 3141 649
rect 3062 631 3064 637
rect 2649 615 2651 621
rect 2944 547 2946 554
rect 2190 514 2192 524
rect 2226 514 2228 524
rect 2234 514 2236 524
rect 2270 514 2272 524
rect 2278 514 2280 524
rect 2321 514 2323 524
rect 2390 520 2392 530
rect 2426 520 2428 530
rect 2434 520 2436 530
rect 2470 520 2472 530
rect 2478 520 2480 530
rect 2521 520 2523 530
rect 2576 529 2578 542
rect 2586 529 2588 542
rect 2618 540 2620 547
rect 3011 543 3013 549
rect 2576 455 2578 468
rect 2586 455 2588 468
rect 2618 466 2620 473
rect 2189 417 2191 427
rect 2225 417 2227 427
rect 2233 417 2235 427
rect 2269 417 2271 427
rect 2277 417 2279 427
rect 2320 417 2322 427
rect 2389 423 2391 433
rect 2425 423 2427 433
rect 2433 423 2435 433
rect 2469 423 2471 433
rect 2477 423 2479 433
rect 2520 423 2522 433
rect 2576 386 2578 399
rect 2586 386 2588 399
rect 2618 397 2620 404
rect 2190 321 2192 331
rect 2226 321 2228 331
rect 2234 321 2236 331
rect 2270 321 2272 331
rect 2278 321 2280 331
rect 2321 321 2323 331
rect 2390 327 2392 337
rect 2426 327 2428 337
rect 2434 327 2436 337
rect 2470 327 2472 337
rect 2478 327 2480 337
rect 2521 327 2523 337
rect 2576 312 2578 325
rect 2586 312 2588 325
rect 2618 323 2620 330
rect 2674 311 2676 535
rect 2681 311 2683 535
rect 2728 312 2730 536
rect 2761 312 2763 536
rect 2792 312 2794 536
rect 2826 313 2828 537
rect 2847 313 2849 537
rect 2869 313 2871 537
rect 2897 314 2899 538
rect 3050 494 3052 506
rect 3060 494 3062 506
rect 3078 494 3080 506
rect 3088 494 3090 506
rect 3165 498 3167 508
rect 3201 498 3203 508
rect 3209 498 3211 508
rect 3245 498 3247 508
rect 3253 498 3255 508
rect 3296 498 3298 508
rect 3011 488 3013 494
rect 2949 471 2951 478
rect 3022 407 3024 413
rect 2952 395 2954 402
rect 3061 358 3063 370
rect 3071 358 3073 370
rect 3089 358 3091 370
rect 3099 358 3101 370
rect 3022 352 3024 358
rect 3178 356 3180 366
rect 3214 356 3216 366
rect 3222 356 3224 366
rect 3258 356 3260 366
rect 3266 356 3268 366
rect 3309 356 3311 366
rect 2941 323 2943 330
rect 3031 273 3033 279
rect 2744 251 2746 261
rect 2787 251 2789 261
rect 2795 251 2797 261
rect 2831 251 2833 261
rect 2839 251 2841 261
rect 2875 251 2877 261
rect 2392 226 2394 236
rect 2428 226 2430 236
rect 2436 226 2438 236
rect 2472 226 2474 236
rect 2480 226 2482 236
rect 2523 226 2525 236
rect 3070 224 3072 236
rect 3080 224 3082 236
rect 3098 224 3100 236
rect 3108 224 3110 236
rect 3188 233 3190 243
rect 3224 233 3226 243
rect 3232 233 3234 243
rect 3268 233 3270 243
rect 3276 233 3278 243
rect 3319 233 3321 243
rect 3031 218 3033 224
rect 3036 124 3038 130
rect 3075 75 3077 87
rect 3085 75 3087 87
rect 3103 75 3105 87
rect 3113 75 3115 87
rect 3193 86 3195 96
rect 3229 86 3231 96
rect 3237 86 3239 96
rect 3273 86 3275 96
rect 3281 86 3283 96
rect 3324 86 3326 96
rect 3036 69 3038 75
<< ptransistor >>
rect 2789 707 2791 719
rect 2649 690 2651 702
rect 2197 647 2199 672
rect 2205 647 2207 672
rect 2235 647 2237 672
rect 2279 647 2281 672
rect 2324 647 2326 672
rect 2392 650 2394 675
rect 2400 650 2402 675
rect 2430 650 2432 675
rect 2474 650 2476 675
rect 2519 650 2521 675
rect 2688 674 2690 698
rect 2698 674 2700 698
rect 2716 668 2718 692
rect 2726 668 2728 692
rect 2828 691 2830 715
rect 2838 691 2840 715
rect 2856 685 2858 709
rect 2866 685 2868 709
rect 2924 707 2926 719
rect 2963 691 2965 715
rect 2973 691 2975 715
rect 2649 635 2651 647
rect 2789 652 2791 664
rect 2991 685 2993 709
rect 3001 685 3003 709
rect 3062 706 3064 718
rect 3101 690 3103 714
rect 3111 690 3113 714
rect 2924 652 2926 664
rect 3129 684 3131 708
rect 3139 684 3141 708
rect 3062 651 3064 663
rect 2782 578 2784 590
rect 2818 579 2820 591
rect 2856 579 2858 591
rect 2194 546 2196 571
rect 2202 546 2204 571
rect 2232 546 2234 571
rect 2276 546 2278 571
rect 2321 546 2323 571
rect 2394 552 2396 577
rect 2402 552 2404 577
rect 2432 552 2434 577
rect 2476 552 2478 577
rect 2521 552 2523 577
rect 2576 565 2578 577
rect 2586 565 2588 577
rect 2618 565 2620 577
rect 2895 578 2897 590
rect 2944 572 2946 584
rect 3011 563 3013 575
rect 3050 547 3052 571
rect 3060 547 3062 571
rect 2576 491 2578 503
rect 2586 491 2588 503
rect 2618 491 2620 503
rect 2193 449 2195 474
rect 2201 449 2203 474
rect 2231 449 2233 474
rect 2275 449 2277 474
rect 2320 449 2322 474
rect 2393 455 2395 480
rect 2401 455 2403 480
rect 2431 455 2433 480
rect 2475 455 2477 480
rect 2520 455 2522 480
rect 2576 422 2578 434
rect 2586 422 2588 434
rect 2618 422 2620 434
rect 2194 353 2196 378
rect 2202 353 2204 378
rect 2232 353 2234 378
rect 2276 353 2278 378
rect 2321 353 2323 378
rect 2394 359 2396 384
rect 2402 359 2404 384
rect 2432 359 2434 384
rect 2476 359 2478 384
rect 2521 359 2523 384
rect 2576 348 2578 360
rect 2586 348 2588 360
rect 2618 348 2620 360
rect 3078 541 3080 565
rect 3088 541 3090 565
rect 3011 508 3013 520
rect 2949 496 2951 508
rect 3169 530 3171 555
rect 3177 530 3179 555
rect 3207 530 3209 555
rect 3251 530 3253 555
rect 3296 530 3298 555
rect 2952 420 2954 432
rect 3022 427 3024 439
rect 3061 411 3063 435
rect 3071 411 3073 435
rect 3089 405 3091 429
rect 3099 405 3101 429
rect 3022 372 3024 384
rect 2941 348 2943 360
rect 3182 388 3184 413
rect 3190 388 3192 413
rect 3220 388 3222 413
rect 3264 388 3266 413
rect 3309 388 3311 413
rect 3031 293 3033 305
rect 2396 258 2398 283
rect 2404 258 2406 283
rect 2434 258 2436 283
rect 2478 258 2480 283
rect 2523 258 2525 283
rect 3070 277 3072 301
rect 3080 277 3082 301
rect 3098 271 3100 295
rect 3108 271 3110 295
rect 3031 238 3033 250
rect 2744 204 2746 229
rect 2789 204 2791 229
rect 2833 204 2835 229
rect 2863 204 2865 229
rect 2871 204 2873 229
rect 3192 265 3194 290
rect 3200 265 3202 290
rect 3230 265 3232 290
rect 3274 265 3276 290
rect 3319 265 3321 290
rect 3036 144 3038 156
rect 3075 128 3077 152
rect 3085 128 3087 152
rect 3103 122 3105 146
rect 3113 122 3115 146
rect 3036 89 3038 101
rect 3197 118 3199 143
rect 3205 118 3207 143
rect 3235 118 3237 143
rect 3279 118 3281 143
rect 3324 118 3326 143
<< ndiffusion >>
rect 2648 670 2649 676
rect 2651 670 2652 676
rect 2788 687 2789 693
rect 2791 687 2792 693
rect 2923 687 2924 693
rect 2926 687 2927 693
rect 2192 615 2193 625
rect 2195 615 2196 625
rect 2228 615 2229 625
rect 2231 615 2232 625
rect 2236 615 2237 625
rect 2239 615 2240 625
rect 2272 615 2273 625
rect 2275 615 2276 625
rect 2280 615 2281 625
rect 2283 615 2284 625
rect 2323 615 2324 625
rect 2326 615 2327 625
rect 2387 618 2388 628
rect 2390 618 2391 628
rect 2423 618 2424 628
rect 2426 618 2427 628
rect 2431 618 2432 628
rect 2434 618 2435 628
rect 2467 618 2468 628
rect 2470 618 2471 628
rect 2475 618 2476 628
rect 2478 618 2479 628
rect 2518 618 2519 628
rect 2521 618 2522 628
rect 3061 686 3062 692
rect 3064 686 3065 692
rect 2827 638 2828 650
rect 2830 638 2838 650
rect 2840 638 2841 650
rect 2855 638 2856 650
rect 2858 638 2866 650
rect 2868 638 2869 650
rect 2962 638 2963 650
rect 2965 638 2973 650
rect 2975 638 2976 650
rect 2990 638 2991 650
rect 2993 638 3001 650
rect 3003 638 3004 650
rect 2687 621 2688 633
rect 2690 621 2698 633
rect 2700 621 2701 633
rect 2715 621 2716 633
rect 2718 621 2726 633
rect 2728 621 2729 633
rect 2788 632 2789 638
rect 2791 632 2792 638
rect 2923 632 2924 638
rect 2926 632 2927 638
rect 3100 637 3101 649
rect 3103 637 3111 649
rect 3113 637 3114 649
rect 3128 637 3129 649
rect 3131 637 3139 649
rect 3141 637 3142 649
rect 3061 631 3062 637
rect 3064 631 3065 637
rect 2648 615 2649 621
rect 2651 615 2652 621
rect 2943 547 2944 554
rect 2946 547 2947 554
rect 2189 514 2190 524
rect 2192 514 2193 524
rect 2225 514 2226 524
rect 2228 514 2229 524
rect 2233 514 2234 524
rect 2236 514 2237 524
rect 2269 514 2270 524
rect 2272 514 2273 524
rect 2277 514 2278 524
rect 2280 514 2281 524
rect 2320 514 2321 524
rect 2323 514 2324 524
rect 2389 520 2390 530
rect 2392 520 2393 530
rect 2425 520 2426 530
rect 2428 520 2429 530
rect 2433 520 2434 530
rect 2436 520 2437 530
rect 2469 520 2470 530
rect 2472 520 2473 530
rect 2477 520 2478 530
rect 2480 520 2481 530
rect 2520 520 2521 530
rect 2523 520 2524 530
rect 2575 529 2576 542
rect 2578 529 2586 542
rect 2588 529 2589 542
rect 2617 540 2618 547
rect 2620 540 2621 547
rect 3010 543 3011 549
rect 3013 543 3014 549
rect 2575 455 2576 468
rect 2578 455 2586 468
rect 2588 455 2589 468
rect 2617 466 2618 473
rect 2620 466 2621 473
rect 2188 417 2189 427
rect 2191 417 2192 427
rect 2224 417 2225 427
rect 2227 417 2228 427
rect 2232 417 2233 427
rect 2235 417 2236 427
rect 2268 417 2269 427
rect 2271 417 2272 427
rect 2276 417 2277 427
rect 2279 417 2280 427
rect 2319 417 2320 427
rect 2322 417 2323 427
rect 2388 423 2389 433
rect 2391 423 2392 433
rect 2424 423 2425 433
rect 2427 423 2428 433
rect 2432 423 2433 433
rect 2435 423 2436 433
rect 2468 423 2469 433
rect 2471 423 2472 433
rect 2476 423 2477 433
rect 2479 423 2480 433
rect 2519 423 2520 433
rect 2522 423 2523 433
rect 2575 386 2576 399
rect 2578 386 2586 399
rect 2588 386 2589 399
rect 2617 397 2618 404
rect 2620 397 2621 404
rect 2189 321 2190 331
rect 2192 321 2193 331
rect 2225 321 2226 331
rect 2228 321 2229 331
rect 2233 321 2234 331
rect 2236 321 2237 331
rect 2269 321 2270 331
rect 2272 321 2273 331
rect 2277 321 2278 331
rect 2280 321 2281 331
rect 2320 321 2321 331
rect 2323 321 2324 331
rect 2389 327 2390 337
rect 2392 327 2393 337
rect 2425 327 2426 337
rect 2428 327 2429 337
rect 2433 327 2434 337
rect 2436 327 2437 337
rect 2469 327 2470 337
rect 2472 327 2473 337
rect 2477 327 2478 337
rect 2480 327 2481 337
rect 2520 327 2521 337
rect 2523 327 2524 337
rect 2575 312 2576 325
rect 2578 312 2586 325
rect 2588 312 2589 325
rect 2617 323 2618 330
rect 2620 323 2621 330
rect 2673 311 2674 535
rect 2676 311 2681 535
rect 2683 311 2684 535
rect 2727 312 2728 536
rect 2730 312 2731 536
rect 2760 312 2761 536
rect 2763 312 2764 536
rect 2791 312 2792 536
rect 2794 312 2795 536
rect 2825 313 2826 537
rect 2828 313 2829 537
rect 2846 313 2847 537
rect 2849 313 2850 537
rect 2868 313 2869 537
rect 2871 313 2872 537
rect 2896 314 2897 538
rect 2899 314 2900 538
rect 3049 494 3050 506
rect 3052 494 3060 506
rect 3062 494 3063 506
rect 3077 494 3078 506
rect 3080 494 3088 506
rect 3090 494 3091 506
rect 3164 498 3165 508
rect 3167 498 3168 508
rect 3200 498 3201 508
rect 3203 498 3204 508
rect 3208 498 3209 508
rect 3211 498 3212 508
rect 3244 498 3245 508
rect 3247 498 3248 508
rect 3252 498 3253 508
rect 3255 498 3256 508
rect 3295 498 3296 508
rect 3298 498 3299 508
rect 3010 488 3011 494
rect 3013 488 3014 494
rect 2948 471 2949 478
rect 2951 471 2952 478
rect 3021 407 3022 413
rect 3024 407 3025 413
rect 2951 395 2952 402
rect 2954 395 2955 402
rect 3060 358 3061 370
rect 3063 358 3071 370
rect 3073 358 3074 370
rect 3088 358 3089 370
rect 3091 358 3099 370
rect 3101 358 3102 370
rect 3021 352 3022 358
rect 3024 352 3025 358
rect 3177 356 3178 366
rect 3180 356 3181 366
rect 3213 356 3214 366
rect 3216 356 3217 366
rect 3221 356 3222 366
rect 3224 356 3225 366
rect 3257 356 3258 366
rect 3260 356 3261 366
rect 3265 356 3266 366
rect 3268 356 3269 366
rect 3308 356 3309 366
rect 3311 356 3312 366
rect 2940 323 2941 330
rect 2943 323 2944 330
rect 3030 273 3031 279
rect 3033 273 3034 279
rect 2743 251 2744 261
rect 2746 251 2747 261
rect 2786 251 2787 261
rect 2789 251 2790 261
rect 2794 251 2795 261
rect 2797 251 2798 261
rect 2830 251 2831 261
rect 2833 251 2834 261
rect 2838 251 2839 261
rect 2841 251 2842 261
rect 2874 251 2875 261
rect 2877 251 2878 261
rect 2391 226 2392 236
rect 2394 226 2395 236
rect 2427 226 2428 236
rect 2430 226 2431 236
rect 2435 226 2436 236
rect 2438 226 2439 236
rect 2471 226 2472 236
rect 2474 226 2475 236
rect 2479 226 2480 236
rect 2482 226 2483 236
rect 2522 226 2523 236
rect 2525 226 2526 236
rect 3069 224 3070 236
rect 3072 224 3080 236
rect 3082 224 3083 236
rect 3097 224 3098 236
rect 3100 224 3108 236
rect 3110 224 3111 236
rect 3187 233 3188 243
rect 3190 233 3191 243
rect 3223 233 3224 243
rect 3226 233 3227 243
rect 3231 233 3232 243
rect 3234 233 3235 243
rect 3267 233 3268 243
rect 3270 233 3271 243
rect 3275 233 3276 243
rect 3278 233 3279 243
rect 3318 233 3319 243
rect 3321 233 3322 243
rect 3030 218 3031 224
rect 3033 218 3034 224
rect 3035 124 3036 130
rect 3038 124 3039 130
rect 3074 75 3075 87
rect 3077 75 3085 87
rect 3087 75 3088 87
rect 3102 75 3103 87
rect 3105 75 3113 87
rect 3115 75 3116 87
rect 3192 86 3193 96
rect 3195 86 3196 96
rect 3228 86 3229 96
rect 3231 86 3232 96
rect 3236 86 3237 96
rect 3239 86 3240 96
rect 3272 86 3273 96
rect 3275 86 3276 96
rect 3280 86 3281 96
rect 3283 86 3284 96
rect 3323 86 3324 96
rect 3326 86 3327 96
rect 3035 69 3036 75
rect 3038 69 3039 75
<< pdiffusion >>
rect 2788 707 2789 719
rect 2791 707 2792 719
rect 2648 690 2649 702
rect 2651 690 2652 702
rect 2196 647 2197 672
rect 2199 647 2200 672
rect 2204 647 2205 672
rect 2207 647 2208 672
rect 2234 647 2235 672
rect 2237 647 2238 672
rect 2278 647 2279 672
rect 2281 647 2282 672
rect 2323 647 2324 672
rect 2326 647 2327 672
rect 2391 650 2392 675
rect 2394 650 2395 675
rect 2399 650 2400 675
rect 2402 650 2403 675
rect 2429 650 2430 675
rect 2432 650 2433 675
rect 2473 650 2474 675
rect 2476 650 2477 675
rect 2518 650 2519 675
rect 2521 650 2522 675
rect 2687 674 2688 698
rect 2690 674 2692 698
rect 2696 674 2698 698
rect 2700 674 2701 698
rect 2715 668 2716 692
rect 2718 668 2720 692
rect 2724 668 2726 692
rect 2728 668 2729 692
rect 2827 691 2828 715
rect 2830 691 2832 715
rect 2836 691 2838 715
rect 2840 691 2841 715
rect 2855 685 2856 709
rect 2858 685 2860 709
rect 2864 685 2866 709
rect 2868 685 2869 709
rect 2923 707 2924 719
rect 2926 707 2927 719
rect 2962 691 2963 715
rect 2965 691 2967 715
rect 2971 691 2973 715
rect 2975 691 2976 715
rect 2648 635 2649 647
rect 2651 635 2652 647
rect 2788 652 2789 664
rect 2791 652 2792 664
rect 2990 685 2991 709
rect 2993 685 2995 709
rect 2999 685 3001 709
rect 3003 685 3004 709
rect 3061 706 3062 718
rect 3064 706 3065 718
rect 3100 690 3101 714
rect 3103 690 3105 714
rect 3109 690 3111 714
rect 3113 690 3114 714
rect 2923 652 2924 664
rect 2926 652 2927 664
rect 3128 684 3129 708
rect 3131 684 3133 708
rect 3137 684 3139 708
rect 3141 684 3142 708
rect 3061 651 3062 663
rect 3064 651 3065 663
rect 2781 578 2782 590
rect 2784 578 2785 590
rect 2817 579 2818 591
rect 2820 579 2821 591
rect 2855 579 2856 591
rect 2858 579 2859 591
rect 2193 546 2194 571
rect 2196 546 2197 571
rect 2201 546 2202 571
rect 2204 546 2205 571
rect 2231 546 2232 571
rect 2234 546 2235 571
rect 2275 546 2276 571
rect 2278 546 2279 571
rect 2320 546 2321 571
rect 2323 546 2324 571
rect 2393 552 2394 577
rect 2396 552 2397 577
rect 2401 552 2402 577
rect 2404 552 2405 577
rect 2431 552 2432 577
rect 2434 552 2435 577
rect 2475 552 2476 577
rect 2478 552 2479 577
rect 2520 552 2521 577
rect 2523 552 2524 577
rect 2575 565 2576 577
rect 2578 565 2580 577
rect 2584 565 2586 577
rect 2588 565 2589 577
rect 2617 565 2618 577
rect 2620 565 2621 577
rect 2894 578 2895 590
rect 2897 578 2898 590
rect 2943 572 2944 584
rect 2946 572 2947 584
rect 3010 563 3011 575
rect 3013 563 3014 575
rect 3049 547 3050 571
rect 3052 547 3054 571
rect 3058 547 3060 571
rect 3062 547 3063 571
rect 2575 491 2576 503
rect 2578 491 2580 503
rect 2584 491 2586 503
rect 2588 491 2589 503
rect 2617 491 2618 503
rect 2620 491 2621 503
rect 2192 449 2193 474
rect 2195 449 2196 474
rect 2200 449 2201 474
rect 2203 449 2204 474
rect 2230 449 2231 474
rect 2233 449 2234 474
rect 2274 449 2275 474
rect 2277 449 2278 474
rect 2319 449 2320 474
rect 2322 449 2323 474
rect 2392 455 2393 480
rect 2395 455 2396 480
rect 2400 455 2401 480
rect 2403 455 2404 480
rect 2430 455 2431 480
rect 2433 455 2434 480
rect 2474 455 2475 480
rect 2477 455 2478 480
rect 2519 455 2520 480
rect 2522 455 2523 480
rect 2575 422 2576 434
rect 2578 422 2580 434
rect 2584 422 2586 434
rect 2588 422 2589 434
rect 2617 422 2618 434
rect 2620 422 2621 434
rect 2193 353 2194 378
rect 2196 353 2197 378
rect 2201 353 2202 378
rect 2204 353 2205 378
rect 2231 353 2232 378
rect 2234 353 2235 378
rect 2275 353 2276 378
rect 2278 353 2279 378
rect 2320 353 2321 378
rect 2323 353 2324 378
rect 2393 359 2394 384
rect 2396 359 2397 384
rect 2401 359 2402 384
rect 2404 359 2405 384
rect 2431 359 2432 384
rect 2434 359 2435 384
rect 2475 359 2476 384
rect 2478 359 2479 384
rect 2520 359 2521 384
rect 2523 359 2524 384
rect 2575 348 2576 360
rect 2578 348 2580 360
rect 2584 348 2586 360
rect 2588 348 2589 360
rect 2617 348 2618 360
rect 2620 348 2621 360
rect 3077 541 3078 565
rect 3080 541 3082 565
rect 3086 541 3088 565
rect 3090 541 3091 565
rect 3010 508 3011 520
rect 3013 508 3014 520
rect 2948 496 2949 508
rect 2951 496 2952 508
rect 3168 530 3169 555
rect 3171 530 3172 555
rect 3176 530 3177 555
rect 3179 530 3180 555
rect 3206 530 3207 555
rect 3209 530 3210 555
rect 3250 530 3251 555
rect 3253 530 3254 555
rect 3295 530 3296 555
rect 3298 530 3299 555
rect 2951 420 2952 432
rect 2954 420 2955 432
rect 3021 427 3022 439
rect 3024 427 3025 439
rect 3060 411 3061 435
rect 3063 411 3065 435
rect 3069 411 3071 435
rect 3073 411 3074 435
rect 3088 405 3089 429
rect 3091 405 3093 429
rect 3097 405 3099 429
rect 3101 405 3102 429
rect 3021 372 3022 384
rect 3024 372 3025 384
rect 2940 348 2941 360
rect 2943 348 2944 360
rect 3181 388 3182 413
rect 3184 388 3185 413
rect 3189 388 3190 413
rect 3192 388 3193 413
rect 3219 388 3220 413
rect 3222 388 3223 413
rect 3263 388 3264 413
rect 3266 388 3267 413
rect 3308 388 3309 413
rect 3311 388 3312 413
rect 3030 293 3031 305
rect 3033 293 3034 305
rect 2395 258 2396 283
rect 2398 258 2399 283
rect 2403 258 2404 283
rect 2406 258 2407 283
rect 2433 258 2434 283
rect 2436 258 2437 283
rect 2477 258 2478 283
rect 2480 258 2481 283
rect 2522 258 2523 283
rect 2525 258 2526 283
rect 3069 277 3070 301
rect 3072 277 3074 301
rect 3078 277 3080 301
rect 3082 277 3083 301
rect 3097 271 3098 295
rect 3100 271 3102 295
rect 3106 271 3108 295
rect 3110 271 3111 295
rect 3030 238 3031 250
rect 3033 238 3034 250
rect 2743 204 2744 229
rect 2746 204 2747 229
rect 2788 204 2789 229
rect 2791 204 2792 229
rect 2832 204 2833 229
rect 2835 204 2836 229
rect 2862 204 2863 229
rect 2865 204 2866 229
rect 2870 204 2871 229
rect 2873 204 2874 229
rect 3191 265 3192 290
rect 3194 265 3195 290
rect 3199 265 3200 290
rect 3202 265 3203 290
rect 3229 265 3230 290
rect 3232 265 3233 290
rect 3273 265 3274 290
rect 3276 265 3277 290
rect 3318 265 3319 290
rect 3321 265 3322 290
rect 3035 144 3036 156
rect 3038 144 3039 156
rect 3074 128 3075 152
rect 3077 128 3079 152
rect 3083 128 3085 152
rect 3087 128 3088 152
rect 3102 122 3103 146
rect 3105 122 3107 146
rect 3111 122 3113 146
rect 3115 122 3116 146
rect 3035 89 3036 101
rect 3038 89 3039 101
rect 3196 118 3197 143
rect 3199 118 3200 143
rect 3204 118 3205 143
rect 3207 118 3208 143
rect 3234 118 3235 143
rect 3237 118 3238 143
rect 3278 118 3279 143
rect 3281 118 3282 143
rect 3323 118 3324 143
rect 3326 118 3327 143
<< ndcontact >>
rect 2644 670 2648 676
rect 2652 670 2656 676
rect 2784 687 2788 693
rect 2792 687 2796 693
rect 2919 687 2923 693
rect 2927 687 2931 693
rect 2188 615 2192 625
rect 2196 615 2200 625
rect 2224 615 2228 625
rect 2232 615 2236 625
rect 2240 615 2244 625
rect 2268 615 2272 625
rect 2276 615 2280 625
rect 2284 615 2288 625
rect 2319 615 2323 625
rect 2327 615 2331 625
rect 2383 618 2387 628
rect 2391 618 2395 628
rect 2419 618 2423 628
rect 2427 618 2431 628
rect 2435 618 2439 628
rect 2463 618 2467 628
rect 2471 618 2475 628
rect 2479 618 2483 628
rect 2514 618 2518 628
rect 2522 618 2526 628
rect 3057 686 3061 692
rect 3065 686 3069 692
rect 2823 638 2827 650
rect 2841 638 2845 650
rect 2851 638 2855 650
rect 2869 638 2873 650
rect 2958 638 2962 650
rect 2976 638 2980 650
rect 2986 638 2990 650
rect 3004 638 3008 650
rect 2683 621 2687 633
rect 2701 621 2705 633
rect 2711 621 2715 633
rect 2729 621 2733 633
rect 2784 632 2788 638
rect 2792 632 2796 638
rect 2919 632 2923 638
rect 2927 632 2931 638
rect 3096 637 3100 649
rect 3114 637 3118 649
rect 3124 637 3128 649
rect 3142 637 3146 649
rect 3057 631 3061 637
rect 3065 631 3069 637
rect 2644 615 2648 621
rect 2652 615 2656 621
rect 2939 547 2943 554
rect 2947 547 2951 554
rect 2185 514 2189 524
rect 2193 514 2197 524
rect 2221 514 2225 524
rect 2229 514 2233 524
rect 2237 514 2241 524
rect 2265 514 2269 524
rect 2273 514 2277 524
rect 2281 514 2285 524
rect 2316 514 2320 524
rect 2324 514 2328 524
rect 2385 520 2389 530
rect 2393 520 2397 530
rect 2421 520 2425 530
rect 2429 520 2433 530
rect 2437 520 2441 530
rect 2465 520 2469 530
rect 2473 520 2477 530
rect 2481 520 2485 530
rect 2516 520 2520 530
rect 2524 520 2528 530
rect 2571 529 2575 542
rect 2589 529 2593 542
rect 2613 540 2617 547
rect 2621 540 2625 547
rect 3006 543 3010 549
rect 3014 543 3018 549
rect 2571 455 2575 468
rect 2589 455 2593 468
rect 2613 466 2617 473
rect 2621 466 2625 473
rect 2184 417 2188 427
rect 2192 417 2196 427
rect 2220 417 2224 427
rect 2228 417 2232 427
rect 2236 417 2240 427
rect 2264 417 2268 427
rect 2272 417 2276 427
rect 2280 417 2284 427
rect 2315 417 2319 427
rect 2323 417 2327 427
rect 2384 423 2388 433
rect 2392 423 2396 433
rect 2420 423 2424 433
rect 2428 423 2432 433
rect 2436 423 2440 433
rect 2464 423 2468 433
rect 2472 423 2476 433
rect 2480 423 2484 433
rect 2515 423 2519 433
rect 2523 423 2527 433
rect 2571 386 2575 399
rect 2589 386 2593 399
rect 2613 397 2617 404
rect 2621 397 2625 404
rect 2185 321 2189 331
rect 2193 321 2197 331
rect 2221 321 2225 331
rect 2229 321 2233 331
rect 2237 321 2241 331
rect 2265 321 2269 331
rect 2273 321 2277 331
rect 2281 321 2285 331
rect 2316 321 2320 331
rect 2324 321 2328 331
rect 2385 327 2389 337
rect 2393 327 2397 337
rect 2421 327 2425 337
rect 2429 327 2433 337
rect 2437 327 2441 337
rect 2465 327 2469 337
rect 2473 327 2477 337
rect 2481 327 2485 337
rect 2516 327 2520 337
rect 2524 327 2528 337
rect 2571 312 2575 325
rect 2589 312 2593 325
rect 2613 323 2617 330
rect 2621 323 2625 330
rect 2669 311 2673 535
rect 2684 311 2689 535
rect 2723 312 2727 536
rect 2731 312 2735 536
rect 2756 312 2760 536
rect 2764 312 2768 536
rect 2787 312 2791 536
rect 2795 312 2799 536
rect 2821 313 2825 537
rect 2829 313 2833 537
rect 2842 313 2846 537
rect 2850 313 2854 537
rect 2864 313 2868 537
rect 2872 313 2876 537
rect 2892 314 2896 538
rect 2900 314 2904 538
rect 3045 494 3049 506
rect 3063 494 3067 506
rect 3073 494 3077 506
rect 3091 494 3095 506
rect 3160 498 3164 508
rect 3168 498 3172 508
rect 3196 498 3200 508
rect 3204 498 3208 508
rect 3212 498 3216 508
rect 3240 498 3244 508
rect 3248 498 3252 508
rect 3256 498 3260 508
rect 3291 498 3295 508
rect 3299 498 3303 508
rect 3006 488 3010 494
rect 3014 488 3018 494
rect 2944 471 2948 478
rect 2952 471 2956 478
rect 3017 407 3021 413
rect 3025 407 3029 413
rect 2947 395 2951 402
rect 2955 395 2959 402
rect 3056 358 3060 370
rect 3074 358 3078 370
rect 3084 358 3088 370
rect 3102 358 3106 370
rect 3017 352 3021 358
rect 3025 352 3029 358
rect 3173 356 3177 366
rect 3181 356 3185 366
rect 3209 356 3213 366
rect 3217 356 3221 366
rect 3225 356 3229 366
rect 3253 356 3257 366
rect 3261 356 3265 366
rect 3269 356 3273 366
rect 3304 356 3308 366
rect 3312 356 3316 366
rect 2936 323 2940 330
rect 2944 323 2948 330
rect 3026 273 3030 279
rect 3034 273 3038 279
rect 2739 251 2743 261
rect 2747 251 2751 261
rect 2782 251 2786 261
rect 2790 251 2794 261
rect 2798 251 2802 261
rect 2826 251 2830 261
rect 2834 251 2838 261
rect 2842 251 2846 261
rect 2870 251 2874 261
rect 2878 251 2882 261
rect 2387 226 2391 236
rect 2395 226 2399 236
rect 2423 226 2427 236
rect 2431 226 2435 236
rect 2439 226 2443 236
rect 2467 226 2471 236
rect 2475 226 2479 236
rect 2483 226 2487 236
rect 2518 226 2522 236
rect 2526 226 2530 236
rect 3065 224 3069 236
rect 3083 224 3087 236
rect 3093 224 3097 236
rect 3111 224 3115 236
rect 3183 233 3187 243
rect 3191 233 3195 243
rect 3219 233 3223 243
rect 3227 233 3231 243
rect 3235 233 3239 243
rect 3263 233 3267 243
rect 3271 233 3275 243
rect 3279 233 3283 243
rect 3314 233 3318 243
rect 3322 233 3326 243
rect 3026 218 3030 224
rect 3034 218 3038 224
rect 3031 124 3035 130
rect 3039 124 3043 130
rect 3070 75 3074 87
rect 3088 75 3092 87
rect 3098 75 3102 87
rect 3116 75 3120 87
rect 3188 86 3192 96
rect 3196 86 3200 96
rect 3224 86 3228 96
rect 3232 86 3236 96
rect 3240 86 3244 96
rect 3268 86 3272 96
rect 3276 86 3280 96
rect 3284 86 3288 96
rect 3319 86 3323 96
rect 3327 86 3331 96
rect 3031 69 3035 75
rect 3039 69 3043 75
<< pdcontact >>
rect 2784 707 2788 719
rect 2792 707 2796 719
rect 2644 690 2648 702
rect 2652 690 2656 702
rect 2192 647 2196 672
rect 2200 647 2204 672
rect 2208 647 2212 672
rect 2230 647 2234 672
rect 2238 647 2242 672
rect 2274 647 2278 672
rect 2282 647 2286 672
rect 2319 647 2323 672
rect 2327 647 2331 672
rect 2387 650 2391 675
rect 2395 650 2399 675
rect 2403 650 2407 675
rect 2425 650 2429 675
rect 2433 650 2437 675
rect 2469 650 2473 675
rect 2477 650 2481 675
rect 2514 650 2518 675
rect 2522 650 2526 675
rect 2683 674 2687 698
rect 2692 674 2696 698
rect 2701 674 2705 698
rect 2711 668 2715 692
rect 2720 668 2724 692
rect 2729 668 2733 692
rect 2823 691 2827 715
rect 2832 691 2836 715
rect 2841 691 2845 715
rect 2851 685 2855 709
rect 2860 685 2864 709
rect 2869 685 2873 709
rect 2919 707 2923 719
rect 2927 707 2931 719
rect 2958 691 2962 715
rect 2967 691 2971 715
rect 2976 691 2980 715
rect 2644 635 2648 647
rect 2652 635 2656 647
rect 2784 652 2788 664
rect 2792 652 2796 664
rect 2986 685 2990 709
rect 2995 685 2999 709
rect 3004 685 3008 709
rect 3057 706 3061 718
rect 3065 706 3069 718
rect 3096 690 3100 714
rect 3105 690 3109 714
rect 3114 690 3118 714
rect 2919 652 2923 664
rect 2927 652 2931 664
rect 3124 684 3128 708
rect 3133 684 3137 708
rect 3142 684 3146 708
rect 3057 651 3061 663
rect 3065 651 3069 663
rect 2777 578 2781 590
rect 2785 578 2789 590
rect 2813 579 2817 591
rect 2821 579 2825 591
rect 2851 579 2855 591
rect 2859 579 2863 591
rect 2189 546 2193 571
rect 2197 546 2201 571
rect 2205 546 2209 571
rect 2227 546 2231 571
rect 2235 546 2239 571
rect 2271 546 2275 571
rect 2279 546 2283 571
rect 2316 546 2320 571
rect 2324 546 2328 571
rect 2389 552 2393 577
rect 2397 552 2401 577
rect 2405 552 2409 577
rect 2427 552 2431 577
rect 2435 552 2439 577
rect 2471 552 2475 577
rect 2479 552 2483 577
rect 2516 552 2520 577
rect 2524 552 2528 577
rect 2571 565 2575 577
rect 2580 565 2584 577
rect 2589 565 2593 577
rect 2613 565 2617 577
rect 2621 565 2625 577
rect 2890 578 2894 590
rect 2898 578 2902 590
rect 2939 572 2943 584
rect 2947 572 2951 584
rect 3006 563 3010 575
rect 3014 563 3018 575
rect 3045 547 3049 571
rect 3054 547 3058 571
rect 3063 547 3067 571
rect 2571 491 2575 503
rect 2580 491 2584 503
rect 2589 491 2593 503
rect 2613 491 2617 503
rect 2621 491 2625 503
rect 2188 449 2192 474
rect 2196 449 2200 474
rect 2204 449 2208 474
rect 2226 449 2230 474
rect 2234 449 2238 474
rect 2270 449 2274 474
rect 2278 449 2282 474
rect 2315 449 2319 474
rect 2323 449 2327 474
rect 2388 455 2392 480
rect 2396 455 2400 480
rect 2404 455 2408 480
rect 2426 455 2430 480
rect 2434 455 2438 480
rect 2470 455 2474 480
rect 2478 455 2482 480
rect 2515 455 2519 480
rect 2523 455 2527 480
rect 2571 422 2575 434
rect 2580 422 2584 434
rect 2589 422 2593 434
rect 2613 422 2617 434
rect 2621 422 2625 434
rect 2189 353 2193 378
rect 2197 353 2201 378
rect 2205 353 2209 378
rect 2227 353 2231 378
rect 2235 353 2239 378
rect 2271 353 2275 378
rect 2279 353 2283 378
rect 2316 353 2320 378
rect 2324 353 2328 378
rect 2389 359 2393 384
rect 2397 359 2401 384
rect 2405 359 2409 384
rect 2427 359 2431 384
rect 2435 359 2439 384
rect 2471 359 2475 384
rect 2479 359 2483 384
rect 2516 359 2520 384
rect 2524 359 2528 384
rect 2571 348 2575 360
rect 2580 348 2584 360
rect 2589 348 2593 360
rect 2613 348 2617 360
rect 2621 348 2625 360
rect 3073 541 3077 565
rect 3082 541 3086 565
rect 3091 541 3095 565
rect 3006 508 3010 520
rect 3014 508 3018 520
rect 2944 496 2948 508
rect 2952 496 2956 508
rect 3164 530 3168 555
rect 3172 530 3176 555
rect 3180 530 3184 555
rect 3202 530 3206 555
rect 3210 530 3214 555
rect 3246 530 3250 555
rect 3254 530 3258 555
rect 3291 530 3295 555
rect 3299 530 3303 555
rect 2947 420 2951 432
rect 2955 420 2959 432
rect 3017 427 3021 439
rect 3025 427 3029 439
rect 3056 411 3060 435
rect 3065 411 3069 435
rect 3074 411 3078 435
rect 3084 405 3088 429
rect 3093 405 3097 429
rect 3102 405 3106 429
rect 3017 372 3021 384
rect 3025 372 3029 384
rect 2936 348 2940 360
rect 2944 348 2948 360
rect 3177 388 3181 413
rect 3185 388 3189 413
rect 3193 388 3197 413
rect 3215 388 3219 413
rect 3223 388 3227 413
rect 3259 388 3263 413
rect 3267 388 3271 413
rect 3304 388 3308 413
rect 3312 388 3316 413
rect 3026 293 3030 305
rect 3034 293 3038 305
rect 2391 258 2395 283
rect 2399 258 2403 283
rect 2407 258 2411 283
rect 2429 258 2433 283
rect 2437 258 2441 283
rect 2473 258 2477 283
rect 2481 258 2485 283
rect 2518 258 2522 283
rect 2526 258 2530 283
rect 3065 277 3069 301
rect 3074 277 3078 301
rect 3083 277 3087 301
rect 3093 271 3097 295
rect 3102 271 3106 295
rect 3111 271 3115 295
rect 3026 238 3030 250
rect 3034 238 3038 250
rect 2739 204 2743 229
rect 2747 204 2751 229
rect 2784 204 2788 229
rect 2792 204 2796 229
rect 2828 204 2832 229
rect 2836 204 2840 229
rect 2858 204 2862 229
rect 2866 204 2870 229
rect 2874 204 2878 229
rect 3187 265 3191 290
rect 3195 265 3199 290
rect 3203 265 3207 290
rect 3225 265 3229 290
rect 3233 265 3237 290
rect 3269 265 3273 290
rect 3277 265 3281 290
rect 3314 265 3318 290
rect 3322 265 3326 290
rect 3031 144 3035 156
rect 3039 144 3043 156
rect 3070 128 3074 152
rect 3079 128 3083 152
rect 3088 128 3092 152
rect 3098 122 3102 146
rect 3107 122 3111 146
rect 3116 122 3120 146
rect 3031 89 3035 101
rect 3039 89 3043 101
rect 3192 118 3196 143
rect 3200 118 3204 143
rect 3208 118 3212 143
rect 3230 118 3234 143
rect 3238 118 3242 143
rect 3274 118 3278 143
rect 3282 118 3286 143
rect 3319 118 3323 143
rect 3327 118 3331 143
<< polysilicon >>
rect 2789 719 2791 722
rect 2924 719 2926 722
rect 2828 715 2830 718
rect 2838 715 2840 718
rect 2649 702 2651 705
rect 2688 698 2690 701
rect 2698 698 2700 701
rect 2392 675 2394 678
rect 2400 675 2402 678
rect 2430 675 2432 678
rect 2474 675 2476 678
rect 2519 675 2521 678
rect 2649 676 2651 690
rect 2197 672 2199 675
rect 2205 672 2207 675
rect 2235 672 2237 675
rect 2279 672 2281 675
rect 2324 672 2326 675
rect 2716 692 2718 695
rect 2726 692 2728 695
rect 2789 693 2791 707
rect 2649 667 2651 670
rect 2688 665 2690 674
rect 2698 664 2700 674
rect 2856 709 2858 712
rect 2866 709 2868 712
rect 2789 684 2791 687
rect 2828 682 2830 691
rect 2838 681 2840 691
rect 3062 718 3064 721
rect 2963 715 2965 718
rect 2973 715 2975 718
rect 2924 693 2926 707
rect 2991 709 2993 712
rect 3001 709 3003 712
rect 2197 640 2199 647
rect 2192 636 2199 640
rect 2193 625 2195 636
rect 2205 628 2207 647
rect 2235 639 2237 647
rect 2279 639 2281 647
rect 2229 637 2237 639
rect 2273 637 2281 639
rect 2229 625 2231 637
rect 2237 625 2239 634
rect 2273 625 2275 637
rect 2281 625 2283 634
rect 2324 625 2326 647
rect 2392 643 2394 650
rect 2387 639 2394 643
rect 2388 628 2390 639
rect 2400 631 2402 650
rect 2430 642 2432 650
rect 2474 642 2476 650
rect 2424 640 2432 642
rect 2468 640 2476 642
rect 2424 628 2426 640
rect 2432 628 2434 637
rect 2468 628 2470 640
rect 2476 628 2478 637
rect 2519 628 2521 650
rect 2649 647 2651 650
rect 2649 621 2651 635
rect 2688 633 2690 660
rect 2698 633 2700 659
rect 2716 657 2718 668
rect 2716 633 2718 653
rect 2726 646 2728 668
rect 2789 664 2791 667
rect 2726 633 2728 642
rect 2789 638 2791 652
rect 2828 650 2830 677
rect 2838 650 2840 676
rect 2856 674 2858 685
rect 2856 650 2858 670
rect 2866 663 2868 685
rect 2924 684 2926 687
rect 2963 682 2965 691
rect 2973 681 2975 691
rect 3101 714 3103 717
rect 3111 714 3113 717
rect 3062 692 3064 706
rect 3129 708 3131 711
rect 3139 708 3141 711
rect 2924 664 2926 667
rect 2866 650 2868 659
rect 2924 638 2926 652
rect 2963 650 2965 677
rect 2973 650 2975 676
rect 2991 674 2993 685
rect 2991 650 2993 670
rect 3001 663 3003 685
rect 3062 683 3064 686
rect 3101 681 3103 690
rect 3111 680 3113 690
rect 3062 663 3064 666
rect 3001 650 3003 659
rect 2828 635 2830 638
rect 2838 635 2840 638
rect 2856 635 2858 638
rect 2866 635 2868 638
rect 2963 635 2965 638
rect 2973 635 2975 638
rect 2991 635 2993 638
rect 3001 635 3003 638
rect 3062 637 3064 651
rect 3101 649 3103 676
rect 3111 649 3113 675
rect 3129 673 3131 684
rect 3129 649 3131 669
rect 3139 662 3141 684
rect 3139 649 3141 658
rect 2789 629 2791 632
rect 2924 629 2926 632
rect 3101 634 3103 637
rect 3111 634 3113 637
rect 3129 634 3131 637
rect 3139 634 3141 637
rect 3062 628 3064 631
rect 2388 615 2390 618
rect 2424 615 2426 618
rect 2432 615 2434 618
rect 2468 615 2470 618
rect 2476 615 2478 618
rect 2519 615 2521 618
rect 2688 618 2690 621
rect 2698 618 2700 621
rect 2716 618 2718 621
rect 2726 618 2728 621
rect 2193 612 2195 615
rect 2229 612 2231 615
rect 2237 612 2239 615
rect 2273 612 2275 615
rect 2281 612 2283 615
rect 2324 612 2326 615
rect 2649 612 2651 615
rect 2782 590 2784 593
rect 2818 591 2820 594
rect 2856 591 2858 594
rect 2394 577 2396 580
rect 2402 577 2404 580
rect 2432 577 2434 580
rect 2476 577 2478 580
rect 2521 577 2523 580
rect 2576 577 2578 580
rect 2586 577 2588 580
rect 2618 577 2620 580
rect 2895 590 2897 593
rect 2194 571 2196 574
rect 2202 571 2204 574
rect 2232 571 2234 574
rect 2276 571 2278 574
rect 2321 571 2323 574
rect 2194 539 2196 546
rect 2189 535 2196 539
rect 2190 524 2192 535
rect 2202 527 2204 546
rect 2232 538 2234 546
rect 2276 538 2278 546
rect 2226 536 2234 538
rect 2270 536 2278 538
rect 2226 524 2228 536
rect 2234 524 2236 533
rect 2270 524 2272 536
rect 2278 524 2280 533
rect 2321 524 2323 546
rect 2394 545 2396 552
rect 2389 541 2396 545
rect 2390 530 2392 541
rect 2402 533 2404 552
rect 2432 544 2434 552
rect 2476 544 2478 552
rect 2426 542 2434 544
rect 2470 542 2478 544
rect 2426 530 2428 542
rect 2434 530 2436 539
rect 2470 530 2472 542
rect 2478 530 2480 539
rect 2521 530 2523 552
rect 2576 542 2578 565
rect 2586 542 2588 565
rect 2618 547 2620 565
rect 2782 563 2784 578
rect 2818 564 2820 579
rect 2856 564 2858 579
rect 2944 584 2946 587
rect 2895 563 2897 578
rect 3011 575 3013 578
rect 2944 554 2946 572
rect 3050 571 3052 574
rect 3060 571 3062 574
rect 3011 549 3013 563
rect 2618 537 2620 540
rect 2674 535 2676 543
rect 2681 535 2683 543
rect 2728 536 2730 543
rect 2761 536 2763 543
rect 2792 536 2794 543
rect 2826 537 2828 544
rect 2847 537 2849 544
rect 2869 537 2871 544
rect 2897 538 2899 545
rect 2944 544 2946 547
rect 3078 565 3080 568
rect 3088 565 3090 568
rect 3011 540 3013 543
rect 3050 538 3052 547
rect 2576 525 2578 529
rect 2586 525 2588 529
rect 2390 517 2392 520
rect 2426 517 2428 520
rect 2434 517 2436 520
rect 2470 517 2472 520
rect 2478 517 2480 520
rect 2521 517 2523 520
rect 2190 511 2192 514
rect 2226 511 2228 514
rect 2234 511 2236 514
rect 2270 511 2272 514
rect 2278 511 2280 514
rect 2321 511 2323 514
rect 2576 503 2578 506
rect 2586 503 2588 506
rect 2618 503 2620 506
rect 2393 480 2395 483
rect 2401 480 2403 483
rect 2431 480 2433 483
rect 2475 480 2477 483
rect 2520 480 2522 483
rect 2193 474 2195 477
rect 2201 474 2203 477
rect 2231 474 2233 477
rect 2275 474 2277 477
rect 2320 474 2322 477
rect 2576 468 2578 491
rect 2586 468 2588 491
rect 2618 473 2620 491
rect 2618 463 2620 466
rect 2193 442 2195 449
rect 2188 438 2195 442
rect 2189 427 2191 438
rect 2201 430 2203 449
rect 2231 441 2233 449
rect 2275 441 2277 449
rect 2225 439 2233 441
rect 2269 439 2277 441
rect 2225 427 2227 439
rect 2233 427 2235 436
rect 2269 427 2271 439
rect 2277 427 2279 436
rect 2320 427 2322 449
rect 2393 448 2395 455
rect 2388 444 2395 448
rect 2389 433 2391 444
rect 2401 436 2403 455
rect 2431 447 2433 455
rect 2475 447 2477 455
rect 2425 445 2433 447
rect 2469 445 2477 447
rect 2425 433 2427 445
rect 2433 433 2435 442
rect 2469 433 2471 445
rect 2477 433 2479 442
rect 2520 433 2522 455
rect 2576 451 2578 455
rect 2586 451 2588 455
rect 2576 434 2578 437
rect 2586 434 2588 437
rect 2618 434 2620 437
rect 2389 420 2391 423
rect 2425 420 2427 423
rect 2433 420 2435 423
rect 2469 420 2471 423
rect 2477 420 2479 423
rect 2520 420 2522 423
rect 2189 414 2191 417
rect 2225 414 2227 417
rect 2233 414 2235 417
rect 2269 414 2271 417
rect 2277 414 2279 417
rect 2320 414 2322 417
rect 2576 399 2578 422
rect 2586 399 2588 422
rect 2618 404 2620 422
rect 2394 384 2396 387
rect 2402 384 2404 387
rect 2432 384 2434 387
rect 2476 384 2478 387
rect 2521 384 2523 387
rect 2618 394 2620 397
rect 2194 378 2196 381
rect 2202 378 2204 381
rect 2232 378 2234 381
rect 2276 378 2278 381
rect 2321 378 2323 381
rect 2576 382 2578 386
rect 2586 382 2588 386
rect 2576 360 2578 363
rect 2586 360 2588 363
rect 2618 360 2620 363
rect 2194 346 2196 353
rect 2189 342 2196 346
rect 2190 331 2192 342
rect 2202 334 2204 353
rect 2232 345 2234 353
rect 2276 345 2278 353
rect 2226 343 2234 345
rect 2270 343 2278 345
rect 2226 331 2228 343
rect 2234 331 2236 340
rect 2270 331 2272 343
rect 2278 331 2280 340
rect 2321 331 2323 353
rect 2394 352 2396 359
rect 2389 348 2396 352
rect 2390 337 2392 348
rect 2402 340 2404 359
rect 2432 351 2434 359
rect 2476 351 2478 359
rect 2426 349 2434 351
rect 2470 349 2478 351
rect 2426 337 2428 349
rect 2434 337 2436 346
rect 2470 337 2472 349
rect 2478 337 2480 346
rect 2521 337 2523 359
rect 2390 324 2392 327
rect 2426 324 2428 327
rect 2434 324 2436 327
rect 2470 324 2472 327
rect 2478 324 2480 327
rect 2521 324 2523 327
rect 2576 325 2578 348
rect 2586 325 2588 348
rect 2618 330 2620 348
rect 2190 318 2192 321
rect 2226 318 2228 321
rect 2234 318 2236 321
rect 2270 318 2272 321
rect 2278 318 2280 321
rect 2321 318 2323 321
rect 2618 320 2620 323
rect 2576 308 2578 312
rect 2586 308 2588 312
rect 3060 537 3062 547
rect 3169 555 3171 558
rect 3177 555 3179 558
rect 3207 555 3209 558
rect 3251 555 3253 558
rect 3296 555 3298 558
rect 3011 520 3013 523
rect 2949 508 2951 511
rect 2949 478 2951 496
rect 3011 494 3013 508
rect 3050 506 3052 533
rect 3060 506 3062 532
rect 3078 530 3080 541
rect 3078 506 3080 526
rect 3088 519 3090 541
rect 3169 523 3171 530
rect 3164 519 3171 523
rect 3088 506 3090 515
rect 3165 508 3167 519
rect 3177 511 3179 530
rect 3207 522 3209 530
rect 3251 522 3253 530
rect 3201 520 3209 522
rect 3245 520 3253 522
rect 3201 508 3203 520
rect 3209 508 3211 517
rect 3245 508 3247 520
rect 3253 508 3255 517
rect 3296 508 3298 530
rect 3165 495 3167 498
rect 3201 495 3203 498
rect 3209 495 3211 498
rect 3245 495 3247 498
rect 3253 495 3255 498
rect 3296 495 3298 498
rect 3050 491 3052 494
rect 3060 491 3062 494
rect 3078 491 3080 494
rect 3088 491 3090 494
rect 3011 485 3013 488
rect 2949 468 2951 471
rect 3022 439 3024 442
rect 2952 432 2954 435
rect 3061 435 3063 438
rect 3071 435 3073 438
rect 2952 402 2954 420
rect 3022 413 3024 427
rect 3089 429 3091 432
rect 3099 429 3101 432
rect 3022 404 3024 407
rect 3061 402 3063 411
rect 3071 401 3073 411
rect 3182 413 3184 416
rect 3190 413 3192 416
rect 3220 413 3222 416
rect 3264 413 3266 416
rect 3309 413 3311 416
rect 2952 392 2954 395
rect 3022 384 3024 387
rect 2941 360 2943 363
rect 3022 358 3024 372
rect 3061 370 3063 397
rect 3071 370 3073 396
rect 3089 394 3091 405
rect 3089 370 3091 390
rect 3099 383 3101 405
rect 3182 381 3184 388
rect 3099 370 3101 379
rect 3177 377 3184 381
rect 3178 366 3180 377
rect 3190 369 3192 388
rect 3220 380 3222 388
rect 3264 380 3266 388
rect 3214 378 3222 380
rect 3258 378 3266 380
rect 3214 366 3216 378
rect 3222 366 3224 375
rect 3258 366 3260 378
rect 3266 366 3268 375
rect 3309 366 3311 388
rect 3061 355 3063 358
rect 3071 355 3073 358
rect 3089 355 3091 358
rect 3099 355 3101 358
rect 3178 353 3180 356
rect 3214 353 3216 356
rect 3222 353 3224 356
rect 3258 353 3260 356
rect 3266 353 3268 356
rect 3309 353 3311 356
rect 3022 349 3024 352
rect 2941 330 2943 348
rect 2941 320 2943 323
rect 2674 308 2676 311
rect 2681 308 2683 311
rect 2728 308 2730 312
rect 2761 308 2763 312
rect 2792 308 2794 312
rect 2826 309 2828 313
rect 2847 309 2849 313
rect 2869 309 2871 313
rect 2897 310 2899 314
rect 3031 305 3033 308
rect 3070 301 3072 304
rect 3080 301 3082 304
rect 2396 283 2398 286
rect 2404 283 2406 286
rect 2434 283 2436 286
rect 2478 283 2480 286
rect 2523 283 2525 286
rect 3031 279 3033 293
rect 3098 295 3100 298
rect 3108 295 3110 298
rect 3031 270 3033 273
rect 3070 268 3072 277
rect 2744 261 2746 264
rect 2787 261 2789 264
rect 2795 261 2797 264
rect 2831 261 2833 264
rect 2839 261 2841 264
rect 2875 261 2877 264
rect 3080 267 3082 277
rect 3192 290 3194 293
rect 3200 290 3202 293
rect 3230 290 3232 293
rect 3274 290 3276 293
rect 3319 290 3321 293
rect 2396 251 2398 258
rect 2391 247 2398 251
rect 2392 236 2394 247
rect 2404 239 2406 258
rect 2434 250 2436 258
rect 2478 250 2480 258
rect 2428 248 2436 250
rect 2472 248 2480 250
rect 2428 236 2430 248
rect 2436 236 2438 245
rect 2472 236 2474 248
rect 2480 236 2482 245
rect 2523 236 2525 258
rect 2744 229 2746 251
rect 2787 242 2789 251
rect 2795 239 2797 251
rect 2831 242 2833 251
rect 2839 239 2841 251
rect 2789 237 2797 239
rect 2833 237 2841 239
rect 2789 229 2791 237
rect 2833 229 2835 237
rect 2863 229 2865 248
rect 2875 240 2877 251
rect 3031 250 3033 253
rect 2871 236 2878 240
rect 2871 229 2873 236
rect 2392 223 2394 226
rect 2428 223 2430 226
rect 2436 223 2438 226
rect 2472 223 2474 226
rect 2480 223 2482 226
rect 2523 223 2525 226
rect 3031 224 3033 238
rect 3070 236 3072 263
rect 3080 236 3082 262
rect 3098 260 3100 271
rect 3098 236 3100 256
rect 3108 249 3110 271
rect 3192 258 3194 265
rect 3187 254 3194 258
rect 3108 236 3110 245
rect 3188 243 3190 254
rect 3200 246 3202 265
rect 3230 257 3232 265
rect 3274 257 3276 265
rect 3224 255 3232 257
rect 3268 255 3276 257
rect 3224 243 3226 255
rect 3232 243 3234 252
rect 3268 243 3270 255
rect 3276 243 3278 252
rect 3319 243 3321 265
rect 3188 230 3190 233
rect 3224 230 3226 233
rect 3232 230 3234 233
rect 3268 230 3270 233
rect 3276 230 3278 233
rect 3319 230 3321 233
rect 3070 221 3072 224
rect 3080 221 3082 224
rect 3098 221 3100 224
rect 3108 221 3110 224
rect 3031 215 3033 218
rect 2744 201 2746 204
rect 2789 201 2791 204
rect 2833 201 2835 204
rect 2863 201 2865 204
rect 2871 201 2873 204
rect 3036 156 3038 159
rect 3075 152 3077 155
rect 3085 152 3087 155
rect 3036 130 3038 144
rect 3103 146 3105 149
rect 3113 146 3115 149
rect 3036 121 3038 124
rect 3075 119 3077 128
rect 3085 118 3087 128
rect 3197 143 3199 146
rect 3205 143 3207 146
rect 3235 143 3237 146
rect 3279 143 3281 146
rect 3324 143 3326 146
rect 3036 101 3038 104
rect 3036 75 3038 89
rect 3075 87 3077 114
rect 3085 87 3087 113
rect 3103 111 3105 122
rect 3103 87 3105 107
rect 3113 100 3115 122
rect 3197 111 3199 118
rect 3192 107 3199 111
rect 3193 96 3195 107
rect 3205 99 3207 118
rect 3235 110 3237 118
rect 3279 110 3281 118
rect 3229 108 3237 110
rect 3273 108 3281 110
rect 3229 96 3231 108
rect 3237 96 3239 105
rect 3273 96 3275 108
rect 3281 96 3283 105
rect 3324 96 3326 118
rect 3113 87 3115 96
rect 3193 83 3195 86
rect 3229 83 3231 86
rect 3237 83 3239 86
rect 3273 83 3275 86
rect 3281 83 3283 86
rect 3324 83 3326 86
rect 3075 72 3077 75
rect 3085 72 3087 75
rect 3103 72 3105 75
rect 3113 72 3115 75
rect 3036 66 3038 69
<< polycontact >>
rect 2645 679 2649 683
rect 2785 696 2789 700
rect 2920 696 2924 700
rect 2188 636 2192 640
rect 2201 628 2205 632
rect 2212 636 2216 640
rect 2224 628 2229 633
rect 2239 628 2243 632
rect 2268 628 2273 633
rect 2320 633 2324 638
rect 2283 628 2287 632
rect 2383 639 2387 643
rect 2396 631 2400 635
rect 2407 639 2411 643
rect 2419 631 2424 636
rect 2434 631 2438 635
rect 2463 631 2468 636
rect 2515 636 2519 641
rect 2478 631 2482 635
rect 2645 624 2649 628
rect 2714 653 2718 657
rect 2725 642 2729 646
rect 2785 641 2789 645
rect 2854 670 2858 674
rect 3058 695 3062 699
rect 2865 659 2869 663
rect 2920 641 2924 645
rect 2989 670 2993 674
rect 3000 659 3004 663
rect 3058 640 3062 644
rect 3127 669 3131 673
rect 3138 658 3142 662
rect 2572 552 2576 556
rect 2185 535 2189 539
rect 2198 527 2202 531
rect 2209 535 2213 539
rect 2221 527 2226 532
rect 2236 527 2240 531
rect 2265 527 2270 532
rect 2317 532 2321 537
rect 2280 527 2284 531
rect 2385 541 2389 545
rect 2398 533 2402 537
rect 2409 541 2413 545
rect 2421 533 2426 538
rect 2436 533 2440 537
rect 2465 533 2470 538
rect 2517 538 2521 543
rect 2480 533 2484 537
rect 2582 545 2586 549
rect 2614 551 2618 555
rect 2778 563 2782 567
rect 2814 564 2818 568
rect 2852 564 2856 568
rect 2891 563 2895 567
rect 2940 558 2944 562
rect 3007 552 3011 556
rect 2670 539 2674 543
rect 2683 539 2687 543
rect 2724 539 2728 543
rect 2757 539 2761 543
rect 2788 539 2792 543
rect 2822 540 2826 544
rect 2843 540 2847 544
rect 2865 540 2869 544
rect 2893 541 2897 545
rect 2572 478 2576 482
rect 2582 471 2586 475
rect 2614 477 2618 481
rect 2184 438 2188 442
rect 2197 430 2201 434
rect 2208 438 2212 442
rect 2220 430 2225 435
rect 2235 430 2239 434
rect 2264 430 2269 435
rect 2316 435 2320 440
rect 2279 430 2283 434
rect 2384 444 2388 448
rect 2397 436 2401 440
rect 2408 444 2412 448
rect 2420 436 2425 441
rect 2435 436 2439 440
rect 2464 436 2469 441
rect 2516 441 2520 446
rect 2479 436 2483 440
rect 2572 409 2576 413
rect 2582 402 2586 406
rect 2614 408 2618 412
rect 2185 342 2189 346
rect 2198 334 2202 338
rect 2209 342 2213 346
rect 2221 334 2226 339
rect 2236 334 2240 338
rect 2265 334 2270 339
rect 2317 339 2321 344
rect 2280 334 2284 338
rect 2385 348 2389 352
rect 2398 340 2402 344
rect 2409 348 2413 352
rect 2421 340 2426 345
rect 2436 340 2440 344
rect 2465 340 2470 345
rect 2517 345 2521 350
rect 2480 340 2484 344
rect 2572 335 2576 339
rect 2582 328 2586 332
rect 2614 334 2618 338
rect 3007 497 3011 501
rect 2945 482 2949 486
rect 3076 526 3080 530
rect 3160 519 3164 523
rect 3087 515 3091 519
rect 3173 511 3177 515
rect 3184 519 3188 523
rect 3196 511 3201 516
rect 3211 511 3215 515
rect 3240 511 3245 516
rect 3292 516 3296 521
rect 3255 511 3259 515
rect 2948 406 2952 410
rect 3018 416 3022 420
rect 3018 361 3022 365
rect 3087 390 3091 394
rect 3098 379 3102 383
rect 3173 377 3177 381
rect 3186 369 3190 373
rect 3197 377 3201 381
rect 3209 369 3214 374
rect 3224 369 3228 373
rect 3253 369 3258 374
rect 3305 374 3309 379
rect 3268 369 3272 373
rect 2937 334 2941 338
rect 3027 282 3031 286
rect 2387 247 2391 251
rect 2400 239 2404 243
rect 2411 247 2415 251
rect 2423 239 2428 244
rect 2438 239 2442 243
rect 2467 239 2472 244
rect 2519 244 2523 249
rect 2482 239 2486 243
rect 2783 244 2787 248
rect 2746 238 2750 243
rect 2797 243 2802 248
rect 2827 244 2831 248
rect 2841 243 2846 248
rect 2854 236 2858 240
rect 2865 244 2869 248
rect 2878 236 2882 240
rect 3027 227 3031 231
rect 3096 256 3100 260
rect 3183 254 3187 258
rect 3107 245 3111 249
rect 3196 246 3200 250
rect 3207 254 3211 258
rect 3219 246 3224 251
rect 3234 246 3238 250
rect 3263 246 3268 251
rect 3315 251 3319 256
rect 3278 246 3282 250
rect 3032 133 3036 137
rect 3032 78 3036 82
rect 3101 107 3105 111
rect 3188 107 3192 111
rect 3112 96 3116 100
rect 3201 99 3205 103
rect 3212 107 3216 111
rect 3224 99 3229 104
rect 3239 99 3243 103
rect 3268 99 3273 104
rect 3320 104 3324 109
rect 3283 99 3287 103
<< metal1 >>
rect 2783 725 2811 728
rect 2918 725 2946 728
rect 2784 719 2787 725
rect 2808 724 2811 725
rect 2808 721 2879 724
rect 2643 708 2671 711
rect 2644 702 2647 708
rect 2668 707 2671 708
rect 2668 704 2739 707
rect 2186 678 2339 682
rect 2381 681 2534 685
rect 2192 672 2196 678
rect 2230 672 2234 678
rect 2274 672 2278 678
rect 2319 672 2323 678
rect 2387 675 2391 681
rect 2425 675 2429 681
rect 2469 675 2473 681
rect 2514 675 2518 681
rect 2627 678 2630 681
rect 2635 679 2645 682
rect 2653 682 2656 690
rect 2683 698 2686 704
rect 2702 698 2705 704
rect 2653 679 2674 682
rect 2653 676 2656 679
rect 2242 647 2255 672
rect 2286 647 2299 672
rect 2437 650 2450 675
rect 2481 650 2494 675
rect 2644 666 2647 670
rect 2638 664 2662 666
rect 2638 663 2656 664
rect 2661 663 2662 664
rect 2671 656 2674 679
rect 2712 698 2732 701
rect 2712 692 2715 698
rect 2729 692 2732 698
rect 2767 695 2770 698
rect 2775 696 2785 699
rect 2793 699 2796 707
rect 2823 715 2826 721
rect 2842 715 2845 721
rect 2919 719 2922 725
rect 2943 724 2946 725
rect 3056 724 3084 727
rect 2943 721 3014 724
rect 2793 696 2814 699
rect 2793 693 2796 696
rect 2693 671 2696 674
rect 2693 668 2711 671
rect 2784 683 2787 687
rect 2778 681 2802 683
rect 2778 680 2796 681
rect 2801 680 2802 681
rect 2811 673 2814 696
rect 2852 715 2872 718
rect 2852 709 2855 715
rect 2869 709 2872 715
rect 2833 688 2836 691
rect 2833 685 2851 688
rect 2902 695 2905 698
rect 2910 696 2920 699
rect 2928 699 2931 707
rect 2958 715 2961 721
rect 2977 715 2980 721
rect 3057 718 3060 724
rect 3081 723 3084 724
rect 3081 720 3152 723
rect 2928 696 2949 699
rect 2928 693 2931 696
rect 2861 678 2864 685
rect 2919 683 2922 687
rect 2913 681 2937 683
rect 2913 680 2931 681
rect 2861 675 2878 678
rect 2783 672 2802 673
rect 2778 670 2802 672
rect 2811 670 2854 673
rect 2721 661 2724 668
rect 2784 664 2787 670
rect 2875 664 2878 675
rect 2936 680 2937 681
rect 2946 673 2949 696
rect 2987 715 3007 718
rect 2987 709 2990 715
rect 3004 709 3007 715
rect 2968 688 2971 691
rect 2968 685 2986 688
rect 3040 694 3043 697
rect 3048 695 3058 698
rect 3066 698 3069 706
rect 3096 714 3099 720
rect 3115 714 3118 720
rect 3066 695 3087 698
rect 3066 692 3069 695
rect 2996 678 2999 685
rect 3057 682 3060 686
rect 3051 680 3075 682
rect 3051 679 3069 680
rect 2996 675 3013 678
rect 2918 672 2937 673
rect 2913 670 2937 672
rect 2946 670 2989 673
rect 2919 664 2922 670
rect 3010 664 3013 675
rect 3074 679 3075 680
rect 3084 672 3087 695
rect 3125 714 3145 717
rect 3125 708 3128 714
rect 3142 708 3145 714
rect 3106 687 3109 690
rect 3106 684 3124 687
rect 3134 677 3137 684
rect 3134 674 3151 677
rect 3056 671 3075 672
rect 3051 669 3075 671
rect 3084 669 3127 672
rect 2721 658 2738 661
rect 2643 655 2662 656
rect 2638 653 2662 655
rect 2671 653 2714 656
rect 2181 636 2188 640
rect 2192 628 2201 632
rect 2208 625 2212 647
rect 2216 636 2217 640
rect 2252 638 2255 647
rect 2296 638 2299 647
rect 2252 633 2264 638
rect 2296 633 2320 638
rect 2327 637 2331 647
rect 2376 639 2383 643
rect 2216 631 2224 633
rect 2221 628 2224 631
rect 2243 628 2244 632
rect 2252 625 2255 633
rect 2260 628 2268 633
rect 2287 628 2288 632
rect 2296 625 2299 633
rect 2327 632 2340 637
rect 2327 625 2331 632
rect 2387 631 2396 635
rect 2403 628 2407 650
rect 2411 639 2412 643
rect 2447 641 2450 650
rect 2491 641 2494 650
rect 2447 636 2459 641
rect 2491 636 2515 641
rect 2522 640 2526 650
rect 2644 647 2647 653
rect 2735 647 2738 658
rect 2840 659 2865 662
rect 2875 660 2887 664
rect 2840 657 2843 659
rect 2411 634 2419 636
rect 2416 631 2419 634
rect 2438 631 2439 635
rect 2447 628 2450 636
rect 2455 631 2463 636
rect 2482 631 2483 635
rect 2491 628 2494 636
rect 2522 635 2542 640
rect 2700 642 2725 645
rect 2735 643 2748 647
rect 2700 640 2703 642
rect 2522 628 2526 635
rect 2200 615 2212 625
rect 2244 615 2255 625
rect 2288 615 2299 625
rect 2395 618 2407 628
rect 2439 618 2450 628
rect 2483 618 2494 628
rect 2188 610 2192 615
rect 2224 610 2228 615
rect 2268 610 2272 615
rect 2319 610 2323 615
rect 2383 613 2387 618
rect 2419 613 2423 618
rect 2463 613 2467 618
rect 2514 613 2518 618
rect 2187 606 2331 610
rect 2382 609 2526 613
rect 2537 597 2542 635
rect 2627 624 2630 627
rect 2635 624 2645 627
rect 2653 627 2656 635
rect 2665 637 2703 640
rect 2735 639 2738 643
rect 2665 627 2668 637
rect 2706 636 2738 639
rect 2706 633 2709 636
rect 2653 624 2668 627
rect 2653 621 2656 624
rect 2705 630 2711 633
rect 2644 611 2647 615
rect 2665 614 2670 617
rect 2683 617 2686 621
rect 2730 617 2733 621
rect 2675 614 2739 617
rect 2665 611 2668 614
rect 2638 608 2668 611
rect 2744 610 2748 643
rect 2767 641 2770 644
rect 2775 641 2785 644
rect 2793 644 2796 652
rect 2805 654 2843 657
rect 2875 656 2878 660
rect 2805 644 2808 654
rect 2846 653 2878 656
rect 2846 650 2849 653
rect 2793 641 2808 644
rect 2793 638 2796 641
rect 2845 647 2851 650
rect 2784 628 2787 632
rect 2805 631 2810 634
rect 2823 634 2826 638
rect 2870 634 2873 638
rect 2815 631 2879 634
rect 2805 628 2808 631
rect 2778 625 2808 628
rect 2883 624 2887 660
rect 2975 659 3000 662
rect 3010 660 3021 664
rect 2975 657 2978 659
rect 2902 641 2905 644
rect 2910 641 2920 644
rect 2928 644 2931 652
rect 2940 654 2978 657
rect 3010 656 3013 660
rect 2940 644 2943 654
rect 2981 653 3013 656
rect 2981 650 2984 653
rect 2928 641 2943 644
rect 2928 638 2931 641
rect 2980 647 2986 650
rect 2919 628 2922 632
rect 2940 631 2945 634
rect 2958 634 2961 638
rect 3005 634 3008 638
rect 2950 631 3014 634
rect 2940 628 2943 631
rect 2913 625 2943 628
rect 2823 621 2887 624
rect 2689 606 2748 610
rect 2754 620 2887 621
rect 3017 620 3021 660
rect 3057 663 3060 669
rect 3148 663 3151 674
rect 3113 658 3138 661
rect 3148 659 3163 663
rect 3113 656 3116 658
rect 3040 640 3043 643
rect 3048 640 3058 643
rect 3066 643 3069 651
rect 3078 653 3116 656
rect 3148 655 3151 659
rect 3078 643 3081 653
rect 3119 652 3151 655
rect 3119 649 3122 652
rect 3066 640 3081 643
rect 3066 637 3069 640
rect 3118 646 3124 649
rect 3057 627 3060 631
rect 3078 630 3083 633
rect 3096 633 3099 637
rect 3143 633 3146 637
rect 3088 630 3152 633
rect 3078 627 3081 630
rect 3051 624 3081 627
rect 3159 623 3163 659
rect 2754 617 2827 620
rect 2537 592 2555 597
rect 2383 583 2536 587
rect 2183 577 2336 581
rect 2389 577 2393 583
rect 2427 577 2431 583
rect 2471 577 2475 583
rect 2516 577 2520 583
rect 2189 571 2193 577
rect 2227 571 2231 577
rect 2271 571 2275 577
rect 2316 571 2320 577
rect 2239 546 2252 571
rect 2283 546 2296 571
rect 2439 552 2452 577
rect 2483 552 2496 577
rect 2550 557 2555 592
rect 2563 583 2634 586
rect 2571 577 2575 583
rect 2589 577 2593 583
rect 2613 577 2616 583
rect 2580 562 2583 565
rect 2580 559 2593 562
rect 2550 556 2563 557
rect 2550 552 2572 556
rect 2590 555 2593 559
rect 2622 555 2625 565
rect 2178 535 2185 539
rect 2189 527 2198 531
rect 2205 524 2209 546
rect 2213 535 2214 539
rect 2249 537 2252 546
rect 2293 537 2296 546
rect 2249 532 2261 537
rect 2293 532 2317 537
rect 2324 536 2328 546
rect 2378 541 2385 545
rect 2213 530 2221 532
rect 2218 527 2221 530
rect 2240 527 2241 531
rect 2249 524 2252 532
rect 2257 527 2265 532
rect 2284 527 2285 531
rect 2293 524 2296 532
rect 2324 531 2337 536
rect 2389 533 2398 537
rect 2324 524 2328 531
rect 2405 530 2409 552
rect 2413 541 2414 545
rect 2449 543 2452 552
rect 2493 543 2496 552
rect 2449 538 2461 543
rect 2493 538 2517 543
rect 2524 542 2528 552
rect 2590 551 2614 555
rect 2622 552 2634 555
rect 2563 545 2582 549
rect 2590 542 2593 551
rect 2622 547 2625 552
rect 2413 536 2421 538
rect 2418 533 2421 536
rect 2440 533 2441 537
rect 2449 530 2452 538
rect 2457 533 2465 538
rect 2484 533 2485 537
rect 2493 530 2496 538
rect 2524 537 2543 542
rect 2524 530 2528 537
rect 2197 514 2209 524
rect 2241 514 2252 524
rect 2285 514 2296 524
rect 2397 520 2409 530
rect 2441 520 2452 530
rect 2485 520 2496 530
rect 2385 515 2389 520
rect 2421 515 2425 520
rect 2465 515 2469 520
rect 2516 515 2520 520
rect 2185 509 2189 514
rect 2221 509 2225 514
rect 2265 509 2269 514
rect 2316 509 2320 514
rect 2384 511 2528 515
rect 2184 505 2328 509
rect 2538 501 2543 537
rect 2689 550 2693 606
rect 2754 603 2758 617
rect 2894 616 3021 620
rect 2831 612 2898 616
rect 2764 608 2835 612
rect 2764 606 2768 608
rect 2708 599 2758 603
rect 2761 602 2768 606
rect 2689 546 2696 550
rect 2692 543 2696 546
rect 2571 523 2574 529
rect 2613 523 2616 540
rect 2667 539 2670 543
rect 2687 539 2696 543
rect 2708 543 2712 599
rect 2761 577 2765 602
rect 2770 596 2798 599
rect 2806 597 2834 600
rect 2844 597 2872 600
rect 2777 590 2780 596
rect 2813 591 2816 597
rect 2851 591 2854 597
rect 2883 596 2911 599
rect 2746 573 2765 577
rect 2746 543 2750 573
rect 2770 563 2778 567
rect 2786 550 2789 578
rect 2806 564 2814 568
rect 2822 557 2825 579
rect 2844 564 2852 568
rect 2822 554 2845 557
rect 2842 550 2845 554
rect 2860 552 2863 579
rect 2890 590 2893 596
rect 2932 590 2964 593
rect 2883 563 2891 567
rect 2899 564 2902 578
rect 2939 584 2942 590
rect 3005 581 3033 584
rect 2786 547 2833 550
rect 2842 547 2854 550
rect 2860 548 2876 552
rect 2899 551 2903 564
rect 2948 562 2951 572
rect 3006 575 3009 581
rect 3030 580 3033 581
rect 3030 577 3101 580
rect 2928 558 2940 562
rect 2948 559 2985 562
rect 2948 554 2951 559
rect 2830 544 2833 547
rect 2708 539 2724 543
rect 2746 539 2757 543
rect 2785 539 2788 543
rect 2795 536 2799 543
rect 2819 540 2822 544
rect 2829 537 2833 544
rect 2840 540 2843 544
rect 2850 537 2854 547
rect 2862 540 2865 544
rect 2872 537 2876 548
rect 2890 541 2893 545
rect 2900 538 2904 551
rect 2563 520 2616 523
rect 2563 509 2634 512
rect 2571 503 2575 509
rect 2589 503 2593 509
rect 2538 496 2551 501
rect 2382 486 2535 490
rect 2182 480 2335 484
rect 2388 480 2392 486
rect 2426 480 2430 486
rect 2470 480 2474 486
rect 2515 480 2519 486
rect 2546 483 2551 496
rect 2613 503 2616 509
rect 2580 488 2583 491
rect 2580 485 2593 488
rect 2546 482 2563 483
rect 2188 474 2192 480
rect 2226 474 2230 480
rect 2270 474 2274 480
rect 2315 474 2319 480
rect 2238 449 2251 474
rect 2282 449 2295 474
rect 2438 455 2451 480
rect 2482 455 2495 480
rect 2546 478 2572 482
rect 2590 481 2593 485
rect 2622 481 2625 491
rect 2590 477 2614 481
rect 2622 478 2634 481
rect 2563 471 2582 475
rect 2590 468 2593 477
rect 2622 473 2625 478
rect 2177 438 2184 442
rect 2188 430 2197 434
rect 2204 427 2208 449
rect 2212 438 2213 442
rect 2248 440 2251 449
rect 2292 440 2295 449
rect 2248 435 2260 440
rect 2292 435 2316 440
rect 2323 439 2327 449
rect 2377 444 2384 448
rect 2212 433 2220 435
rect 2217 430 2220 433
rect 2239 430 2240 434
rect 2248 427 2251 435
rect 2256 430 2264 435
rect 2283 430 2284 434
rect 2292 427 2295 435
rect 2323 434 2336 439
rect 2388 436 2397 440
rect 2323 427 2327 434
rect 2404 433 2408 455
rect 2412 444 2413 448
rect 2448 446 2451 455
rect 2492 446 2495 455
rect 2448 441 2460 446
rect 2492 441 2516 446
rect 2523 445 2527 455
rect 2571 449 2574 455
rect 2613 449 2616 466
rect 2563 446 2616 449
rect 2412 439 2420 441
rect 2417 436 2420 439
rect 2439 436 2440 440
rect 2448 433 2451 441
rect 2456 436 2464 441
rect 2483 436 2484 440
rect 2492 433 2495 441
rect 2523 440 2554 445
rect 2563 440 2634 443
rect 2523 433 2527 440
rect 2196 417 2208 427
rect 2240 417 2251 427
rect 2284 417 2295 427
rect 2396 423 2408 433
rect 2440 423 2451 433
rect 2484 423 2495 433
rect 2384 418 2388 423
rect 2420 418 2424 423
rect 2464 418 2468 423
rect 2515 418 2519 423
rect 2184 412 2188 417
rect 2220 412 2224 417
rect 2264 412 2268 417
rect 2315 412 2319 417
rect 2383 414 2527 418
rect 2549 413 2554 440
rect 2571 434 2575 440
rect 2589 434 2593 440
rect 2613 434 2616 440
rect 2580 419 2583 422
rect 2580 416 2593 419
rect 2183 408 2327 412
rect 2549 409 2572 413
rect 2590 412 2593 416
rect 2622 412 2625 422
rect 2590 408 2614 412
rect 2622 409 2634 412
rect 2563 402 2582 406
rect 2590 399 2593 408
rect 2622 404 2625 409
rect 2383 390 2536 394
rect 2183 384 2336 388
rect 2389 384 2393 390
rect 2427 384 2431 390
rect 2471 384 2475 390
rect 2516 384 2520 390
rect 2189 378 2193 384
rect 2227 378 2231 384
rect 2271 378 2275 384
rect 2316 378 2320 384
rect 2239 353 2252 378
rect 2283 353 2296 378
rect 2439 359 2452 384
rect 2483 359 2496 384
rect 2571 380 2574 386
rect 2613 380 2616 397
rect 2563 377 2616 380
rect 2563 366 2634 369
rect 2178 342 2185 346
rect 2189 334 2198 338
rect 2205 331 2209 353
rect 2213 342 2214 346
rect 2249 344 2252 353
rect 2293 344 2296 353
rect 2249 339 2261 344
rect 2293 339 2317 344
rect 2324 343 2328 353
rect 2378 348 2385 352
rect 2213 337 2221 339
rect 2218 334 2221 337
rect 2240 334 2241 338
rect 2249 331 2252 339
rect 2257 334 2265 339
rect 2284 334 2285 338
rect 2293 331 2296 339
rect 2324 338 2337 343
rect 2389 340 2398 344
rect 2324 331 2328 338
rect 2405 337 2409 359
rect 2413 348 2414 352
rect 2449 350 2452 359
rect 2493 350 2496 359
rect 2449 345 2461 350
rect 2493 345 2517 350
rect 2524 349 2528 359
rect 2571 360 2575 366
rect 2589 360 2593 366
rect 2413 343 2421 345
rect 2418 340 2421 343
rect 2440 340 2441 344
rect 2449 337 2452 345
rect 2457 340 2465 345
rect 2484 340 2485 344
rect 2493 337 2496 345
rect 2524 344 2554 349
rect 2613 360 2616 366
rect 2524 337 2528 344
rect 2197 321 2209 331
rect 2241 321 2252 331
rect 2285 321 2296 331
rect 2397 327 2409 337
rect 2441 327 2452 337
rect 2485 327 2496 337
rect 2549 339 2554 344
rect 2580 345 2583 348
rect 2580 342 2593 345
rect 2549 335 2572 339
rect 2590 338 2593 342
rect 2622 338 2625 348
rect 2590 334 2614 338
rect 2622 335 2634 338
rect 2563 328 2582 332
rect 2385 322 2389 327
rect 2421 322 2425 327
rect 2465 322 2469 327
rect 2516 322 2520 327
rect 2590 325 2593 334
rect 2622 330 2625 335
rect 2185 316 2189 321
rect 2221 316 2225 321
rect 2265 316 2269 321
rect 2316 316 2320 321
rect 2384 318 2528 322
rect 2184 312 2328 316
rect 2571 306 2574 312
rect 2613 306 2616 323
rect 2563 303 2616 306
rect 2669 302 2673 311
rect 2684 310 2689 311
rect 2723 310 2727 312
rect 2684 305 2727 310
rect 2731 310 2735 312
rect 2756 310 2760 312
rect 2731 305 2760 310
rect 2764 310 2768 312
rect 2939 530 2942 547
rect 2928 527 2942 530
rect 2933 514 2965 517
rect 2944 508 2947 514
rect 2953 486 2956 496
rect 2933 482 2945 486
rect 2953 483 2979 486
rect 2953 478 2956 483
rect 2944 454 2947 471
rect 2933 451 2947 454
rect 2936 438 2968 441
rect 2947 432 2950 438
rect 2956 410 2959 420
rect 2936 406 2948 410
rect 2956 407 2968 410
rect 2956 402 2959 407
rect 2947 378 2950 395
rect 2965 388 2968 407
rect 2965 385 2972 388
rect 2936 375 2950 378
rect 2925 366 2957 369
rect 2936 360 2939 366
rect 2945 338 2948 348
rect 2925 334 2937 338
rect 2945 335 2962 338
rect 2945 330 2948 335
rect 2787 310 2791 312
rect 2764 305 2791 310
rect 2821 308 2825 313
rect 2842 308 2846 313
rect 2864 308 2868 313
rect 2892 308 2896 314
rect 2821 305 2896 308
rect 2936 306 2939 323
rect 2925 303 2939 306
rect 2664 298 2682 302
rect 2385 289 2538 293
rect 2391 283 2395 289
rect 2429 283 2433 289
rect 2473 283 2477 289
rect 2518 283 2522 289
rect 2441 258 2454 283
rect 2485 258 2498 283
rect 2739 266 2883 270
rect 2747 261 2751 266
rect 2798 261 2802 266
rect 2842 261 2846 266
rect 2878 261 2882 266
rect 2380 247 2387 251
rect 2391 239 2400 243
rect 2407 236 2411 258
rect 2415 247 2416 251
rect 2451 249 2454 258
rect 2495 249 2498 258
rect 2451 244 2463 249
rect 2495 244 2519 249
rect 2526 248 2530 258
rect 2771 251 2782 261
rect 2815 251 2826 261
rect 2858 251 2870 261
rect 2415 242 2423 244
rect 2420 239 2423 242
rect 2442 239 2443 243
rect 2451 236 2454 244
rect 2459 239 2467 244
rect 2486 239 2487 243
rect 2495 236 2498 244
rect 2526 243 2539 248
rect 2739 244 2743 251
rect 2526 236 2530 243
rect 2730 239 2743 244
rect 2771 243 2774 251
rect 2782 244 2783 248
rect 2802 243 2810 248
rect 2815 243 2818 251
rect 2826 244 2827 248
rect 2846 245 2849 248
rect 2846 243 2854 245
rect 2399 226 2411 236
rect 2443 226 2454 236
rect 2487 226 2498 236
rect 2739 229 2743 239
rect 2750 238 2774 243
rect 2806 238 2818 243
rect 2771 229 2774 238
rect 2815 229 2818 238
rect 2853 236 2854 240
rect 2858 229 2862 251
rect 2869 244 2878 248
rect 2959 243 2962 335
rect 2969 334 2972 385
rect 2976 342 2979 483
rect 2982 364 2985 559
rect 2989 551 2992 554
rect 2997 552 3007 555
rect 3015 555 3018 563
rect 3045 571 3048 577
rect 3064 571 3067 577
rect 3015 552 3036 555
rect 3015 549 3018 552
rect 3006 539 3009 543
rect 3000 537 3024 539
rect 3000 536 3018 537
rect 3023 536 3024 537
rect 3033 529 3036 552
rect 3074 571 3094 574
rect 3074 565 3077 571
rect 3091 565 3094 571
rect 3055 544 3058 547
rect 3055 541 3073 544
rect 3158 561 3311 565
rect 3164 555 3168 561
rect 3202 555 3206 561
rect 3246 555 3250 561
rect 3291 555 3295 561
rect 3083 534 3086 541
rect 3083 531 3100 534
rect 3005 528 3024 529
rect 3000 526 3024 528
rect 3033 526 3076 529
rect 3006 520 3009 526
rect 3097 520 3100 531
rect 3214 530 3227 555
rect 3258 530 3271 555
rect 3124 520 3160 523
rect 3097 519 3160 520
rect 3062 515 3087 518
rect 3097 516 3128 519
rect 3062 513 3065 515
rect 2989 497 2992 500
rect 2997 497 3007 500
rect 3015 500 3018 508
rect 3027 510 3065 513
rect 3097 512 3100 516
rect 3027 500 3030 510
rect 3068 509 3100 512
rect 3164 511 3173 515
rect 3068 506 3071 509
rect 3180 508 3184 530
rect 3188 519 3189 523
rect 3224 521 3227 530
rect 3268 521 3271 530
rect 3224 516 3236 521
rect 3268 516 3292 521
rect 3299 520 3303 530
rect 3188 514 3196 516
rect 3193 511 3196 514
rect 3215 511 3216 515
rect 3224 508 3227 516
rect 3232 511 3240 516
rect 3259 511 3260 515
rect 3268 508 3271 516
rect 3299 515 3312 520
rect 3299 508 3303 515
rect 3015 497 3030 500
rect 3015 494 3018 497
rect 3067 503 3073 506
rect 3006 484 3009 488
rect 3027 487 3032 490
rect 3045 490 3048 494
rect 3092 490 3095 494
rect 3172 498 3184 508
rect 3216 498 3227 508
rect 3260 498 3271 508
rect 3160 493 3164 498
rect 3196 493 3200 498
rect 3240 493 3244 498
rect 3291 493 3295 498
rect 3037 487 3101 490
rect 3159 489 3303 493
rect 3027 484 3030 487
rect 3000 481 3030 484
rect 3016 445 3044 448
rect 3017 439 3020 445
rect 3041 444 3044 445
rect 3041 441 3112 444
rect 3000 415 3003 418
rect 3008 416 3018 419
rect 3026 419 3029 427
rect 3056 435 3059 441
rect 3075 435 3078 441
rect 3026 416 3047 419
rect 3026 413 3029 416
rect 3017 403 3020 407
rect 3011 401 3035 403
rect 3011 400 3029 401
rect 3034 400 3035 401
rect 3044 393 3047 416
rect 3085 435 3105 438
rect 3085 429 3088 435
rect 3102 429 3105 435
rect 3066 408 3069 411
rect 3066 405 3084 408
rect 3171 419 3324 423
rect 3177 413 3181 419
rect 3215 413 3219 419
rect 3259 413 3263 419
rect 3304 413 3308 419
rect 3094 398 3097 405
rect 3094 395 3111 398
rect 3016 392 3035 393
rect 3011 390 3035 392
rect 3044 390 3087 393
rect 3017 384 3020 390
rect 3108 384 3111 395
rect 3227 388 3240 413
rect 3271 388 3284 413
rect 3073 379 3098 382
rect 3108 381 3164 384
rect 3108 380 3173 381
rect 3073 377 3076 379
rect 2982 361 3003 364
rect 3008 361 3018 364
rect 3026 364 3029 372
rect 3038 374 3076 377
rect 3108 376 3111 380
rect 3160 377 3173 380
rect 3038 364 3041 374
rect 3079 373 3111 376
rect 3079 370 3082 373
rect 3026 361 3041 364
rect 3026 358 3029 361
rect 3078 367 3084 370
rect 3177 369 3186 373
rect 3193 366 3197 388
rect 3201 377 3202 381
rect 3237 379 3240 388
rect 3281 379 3284 388
rect 3237 374 3249 379
rect 3281 374 3305 379
rect 3312 378 3316 388
rect 3201 372 3209 374
rect 3206 369 3209 372
rect 3228 369 3229 373
rect 3237 366 3240 374
rect 3245 369 3253 374
rect 3272 369 3273 373
rect 3281 366 3284 374
rect 3312 373 3325 378
rect 3312 366 3316 373
rect 3017 348 3020 352
rect 3038 351 3043 354
rect 3056 354 3059 358
rect 3103 354 3106 358
rect 3185 356 3197 366
rect 3229 356 3240 366
rect 3273 356 3284 366
rect 3048 351 3112 354
rect 3173 351 3177 356
rect 3209 351 3213 356
rect 3253 351 3257 356
rect 3304 351 3308 356
rect 3038 348 3041 351
rect 3011 345 3041 348
rect 3172 347 3316 351
rect 2976 339 3005 342
rect 2969 331 2995 334
rect 2911 240 2962 243
rect 2882 236 2915 240
rect 2387 221 2391 226
rect 2423 221 2427 226
rect 2467 221 2471 226
rect 2518 221 2522 226
rect 2386 217 2530 221
rect 2771 204 2784 229
rect 2815 204 2828 229
rect 2747 198 2751 204
rect 2792 198 2796 204
rect 2836 198 2840 204
rect 2874 198 2878 204
rect 2731 194 2884 198
rect 2992 81 2995 331
rect 3002 230 3005 339
rect 3025 311 3053 314
rect 3026 305 3029 311
rect 3050 310 3053 311
rect 3050 307 3121 310
rect 3009 281 3012 284
rect 3017 282 3027 285
rect 3035 285 3038 293
rect 3065 301 3068 307
rect 3084 301 3087 307
rect 3035 282 3056 285
rect 3035 279 3038 282
rect 3026 269 3029 273
rect 3020 267 3044 269
rect 3020 266 3038 267
rect 3043 266 3044 267
rect 3053 259 3056 282
rect 3094 301 3114 304
rect 3094 295 3097 301
rect 3111 295 3114 301
rect 3181 296 3334 300
rect 3075 274 3078 277
rect 3075 271 3093 274
rect 3187 290 3191 296
rect 3225 290 3229 296
rect 3269 290 3273 296
rect 3314 290 3318 296
rect 3103 264 3106 271
rect 3237 265 3250 290
rect 3281 265 3294 290
rect 3103 261 3120 264
rect 3025 258 3044 259
rect 3020 256 3044 258
rect 3053 256 3096 259
rect 3026 250 3029 256
rect 3117 250 3120 261
rect 3151 254 3183 258
rect 3151 250 3155 254
rect 3082 245 3107 248
rect 3117 246 3155 250
rect 3187 246 3196 250
rect 3082 243 3085 245
rect 3002 227 3012 230
rect 3017 227 3027 230
rect 3035 230 3038 238
rect 3047 240 3085 243
rect 3117 242 3120 246
rect 3203 243 3207 265
rect 3211 254 3212 258
rect 3247 256 3250 265
rect 3291 256 3294 265
rect 3247 251 3259 256
rect 3291 251 3315 256
rect 3322 255 3326 265
rect 3211 249 3219 251
rect 3216 246 3219 249
rect 3238 246 3239 250
rect 3247 243 3250 251
rect 3255 246 3263 251
rect 3282 246 3283 250
rect 3291 243 3294 251
rect 3322 250 3335 255
rect 3322 243 3326 250
rect 3047 230 3050 240
rect 3088 239 3120 242
rect 3088 236 3091 239
rect 3035 227 3050 230
rect 3035 224 3038 227
rect 3087 233 3093 236
rect 3195 233 3207 243
rect 3239 233 3250 243
rect 3283 233 3294 243
rect 3183 228 3187 233
rect 3219 228 3223 233
rect 3263 228 3267 233
rect 3314 228 3318 233
rect 3182 224 3326 228
rect 3026 214 3029 218
rect 3047 217 3052 220
rect 3065 220 3068 224
rect 3112 220 3115 224
rect 3057 217 3121 220
rect 3047 214 3050 217
rect 3020 211 3050 214
rect 3030 162 3058 165
rect 3031 156 3034 162
rect 3055 161 3058 162
rect 3055 158 3126 161
rect 3014 132 3017 135
rect 3022 133 3032 136
rect 3040 136 3043 144
rect 3070 152 3073 158
rect 3089 152 3092 158
rect 3040 133 3061 136
rect 3040 130 3043 133
rect 3031 120 3034 124
rect 3025 118 3049 120
rect 3025 117 3043 118
rect 3048 117 3049 118
rect 3058 110 3061 133
rect 3099 152 3119 155
rect 3099 146 3102 152
rect 3116 146 3119 152
rect 3186 149 3339 153
rect 3080 125 3083 128
rect 3080 122 3098 125
rect 3192 143 3196 149
rect 3230 143 3234 149
rect 3274 143 3278 149
rect 3319 143 3323 149
rect 3108 115 3111 122
rect 3242 118 3255 143
rect 3286 118 3299 143
rect 3108 112 3125 115
rect 3030 109 3049 110
rect 3025 107 3049 109
rect 3058 107 3101 110
rect 3031 101 3034 107
rect 3122 101 3125 112
rect 3151 107 3188 111
rect 3151 101 3155 107
rect 3087 96 3112 99
rect 3122 97 3155 101
rect 3192 99 3201 103
rect 3087 94 3090 96
rect 2992 78 3017 81
rect 3022 78 3032 81
rect 3040 81 3043 89
rect 3052 91 3090 94
rect 3122 93 3125 97
rect 3208 96 3212 118
rect 3216 107 3217 111
rect 3252 109 3255 118
rect 3296 109 3299 118
rect 3252 104 3264 109
rect 3296 104 3320 109
rect 3327 108 3331 118
rect 3216 102 3224 104
rect 3221 99 3224 102
rect 3243 99 3244 103
rect 3252 96 3255 104
rect 3260 99 3268 104
rect 3287 99 3288 103
rect 3296 96 3299 104
rect 3327 103 3340 108
rect 3327 96 3331 103
rect 3052 81 3055 91
rect 3093 90 3125 93
rect 3093 87 3096 90
rect 3040 78 3055 81
rect 3040 75 3043 78
rect 3092 84 3098 87
rect 3200 86 3212 96
rect 3244 86 3255 96
rect 3288 86 3299 96
rect 3188 81 3192 86
rect 3224 81 3228 86
rect 3268 81 3272 86
rect 3319 81 3323 86
rect 3187 77 3331 81
rect 3031 65 3034 69
rect 3052 68 3057 71
rect 3070 71 3073 75
rect 3117 71 3120 75
rect 3062 68 3126 71
rect 3052 65 3055 68
rect 3025 62 3055 65
<< m2contact >>
rect 2630 677 2635 682
rect 2770 694 2775 699
rect 2905 694 2910 699
rect 3043 693 3048 698
rect 2187 628 2192 633
rect 2217 636 2222 641
rect 2216 626 2221 631
rect 2244 628 2249 633
rect 2288 628 2293 633
rect 2382 631 2387 636
rect 2412 639 2417 644
rect 2411 629 2416 634
rect 2439 631 2444 636
rect 2483 631 2488 636
rect 2630 623 2635 628
rect 2770 640 2775 645
rect 2905 640 2910 645
rect 3043 639 3048 644
rect 2184 527 2189 532
rect 2214 535 2219 540
rect 2213 525 2218 530
rect 2241 527 2246 532
rect 2285 527 2290 532
rect 2384 533 2389 538
rect 2414 541 2419 546
rect 2413 531 2418 536
rect 2441 533 2446 538
rect 2485 533 2490 538
rect 2789 559 2794 564
rect 2845 550 2850 555
rect 2923 558 2928 563
rect 2876 541 2881 546
rect 2183 430 2188 435
rect 2213 438 2218 443
rect 2212 428 2217 433
rect 2240 430 2245 435
rect 2284 430 2289 435
rect 2383 436 2388 441
rect 2413 444 2418 449
rect 2412 434 2417 439
rect 2440 436 2445 441
rect 2484 436 2489 441
rect 2184 334 2189 339
rect 2214 342 2219 347
rect 2213 332 2218 337
rect 2241 334 2246 339
rect 2285 334 2290 339
rect 2384 340 2389 345
rect 2414 348 2419 353
rect 2413 338 2418 343
rect 2441 340 2446 345
rect 2485 340 2490 345
rect 2928 482 2933 487
rect 2931 406 2936 411
rect 2386 239 2391 244
rect 2416 247 2421 252
rect 2415 237 2420 242
rect 2443 239 2448 244
rect 2487 239 2492 244
rect 2777 243 2782 248
rect 2821 243 2826 248
rect 2849 245 2854 250
rect 2848 235 2853 240
rect 2878 243 2883 248
rect 2992 550 2997 555
rect 2992 496 2997 501
rect 3159 511 3164 516
rect 3189 519 3194 524
rect 3188 509 3193 514
rect 3216 511 3221 516
rect 3260 511 3265 516
rect 3003 414 3008 419
rect 3003 360 3008 365
rect 3172 369 3177 374
rect 3202 377 3207 382
rect 3201 367 3206 372
rect 3229 369 3234 374
rect 3273 369 3278 374
rect 3012 280 3017 285
rect 3182 246 3187 251
rect 3012 226 3017 231
rect 3212 254 3217 259
rect 3211 244 3216 249
rect 3239 246 3244 251
rect 3283 246 3288 251
rect 3017 131 3022 136
rect 3187 99 3192 104
rect 3017 77 3022 82
rect 3217 107 3222 112
rect 3216 97 3221 102
rect 3244 99 3249 104
rect 3288 99 3293 104
<< pm12contact >>
rect 2826 677 2831 682
rect 2835 676 2840 681
rect 2686 660 2691 665
rect 2695 659 2700 664
rect 2961 677 2966 682
rect 2970 676 2975 681
rect 3099 676 3104 681
rect 3108 675 3113 680
rect 3048 533 3053 538
rect 3057 532 3062 537
rect 3059 397 3064 402
rect 3068 396 3073 401
rect 3068 263 3073 268
rect 3077 262 3082 267
rect 3073 114 3078 119
rect 3082 113 3087 118
<< metal2 >>
rect 2412 689 2443 692
rect 2217 686 2248 689
rect 2217 641 2221 686
rect 2244 633 2248 686
rect 2412 644 2416 689
rect 2166 628 2187 632
rect 2178 604 2184 628
rect 2439 636 2443 689
rect 2771 688 2774 694
rect 2906 688 2909 694
rect 2771 685 2808 688
rect 2906 685 2943 688
rect 2805 682 2808 685
rect 2940 682 2943 685
rect 3044 687 3047 693
rect 3044 684 3081 687
rect 2631 671 2634 677
rect 2805 679 2826 682
rect 2631 668 2668 671
rect 2665 665 2668 668
rect 2835 666 2838 676
rect 2940 679 2961 682
rect 3078 681 3081 684
rect 2970 666 2973 676
rect 3078 678 3099 681
rect 2665 662 2686 665
rect 2772 663 2838 666
rect 2907 663 2973 666
rect 3108 665 3111 675
rect 2695 649 2698 659
rect 2632 646 2698 649
rect 2361 631 2382 635
rect 2217 604 2221 626
rect 2288 604 2293 628
rect 2373 607 2379 631
rect 2412 607 2416 629
rect 2483 607 2488 631
rect 2632 628 2635 646
rect 2772 645 2775 663
rect 2907 645 2910 663
rect 3045 662 3111 665
rect 3045 644 3048 662
rect 2373 604 2492 607
rect 2178 601 2297 604
rect 2414 591 2445 594
rect 2214 585 2245 588
rect 2214 540 2218 585
rect 2241 532 2245 585
rect 2414 546 2418 591
rect 2441 538 2445 591
rect 3189 569 3220 572
rect 2794 559 2923 563
rect 2850 550 2927 554
rect 2876 538 2881 541
rect 2163 527 2184 531
rect 2175 503 2181 527
rect 2363 533 2384 537
rect 2214 503 2218 525
rect 2285 503 2290 527
rect 2375 509 2381 533
rect 2414 509 2418 531
rect 2485 509 2490 533
rect 2375 506 2494 509
rect 2175 500 2294 503
rect 2413 494 2444 497
rect 2213 488 2244 491
rect 2213 443 2217 488
rect 2240 435 2244 488
rect 2413 449 2417 494
rect 2440 441 2444 494
rect 2162 430 2183 434
rect 2174 406 2180 430
rect 2362 436 2383 440
rect 2213 406 2217 428
rect 2284 406 2289 430
rect 2374 412 2380 436
rect 2413 412 2417 434
rect 2484 412 2489 436
rect 2374 409 2493 412
rect 2174 403 2293 406
rect 2877 406 2880 538
rect 2923 489 2927 550
rect 2993 544 2996 550
rect 2993 541 3030 544
rect 3027 538 3030 541
rect 3027 535 3048 538
rect 3057 522 3060 532
rect 2994 519 3060 522
rect 3189 524 3193 569
rect 2994 501 2997 519
rect 3216 516 3220 569
rect 3138 511 3159 515
rect 2923 486 2928 489
rect 3150 487 3156 511
rect 3189 487 3193 509
rect 3260 487 3265 511
rect 2925 482 2928 486
rect 3150 484 3269 487
rect 3202 427 3233 430
rect 2927 406 2931 411
rect 3004 408 3007 414
rect 2877 403 2931 406
rect 3004 405 3041 408
rect 3038 402 3041 405
rect 2414 398 2445 401
rect 2214 392 2245 395
rect 2214 347 2218 392
rect 2241 339 2245 392
rect 2414 353 2418 398
rect 2441 345 2445 398
rect 3038 399 3059 402
rect 3068 386 3071 396
rect 3005 383 3071 386
rect 3005 365 3008 383
rect 3202 382 3206 427
rect 3229 374 3233 427
rect 3037 368 3040 371
rect 3151 369 3172 373
rect 3163 345 3169 369
rect 3202 345 3206 367
rect 3273 345 3278 369
rect 2163 334 2184 338
rect 2175 310 2181 334
rect 2363 340 2384 344
rect 2214 310 2218 332
rect 2285 310 2290 334
rect 2375 316 2381 340
rect 3163 342 3282 345
rect 2414 316 2418 338
rect 2485 316 2490 340
rect 2375 313 2494 316
rect 2175 307 2294 310
rect 3212 304 3243 307
rect 2416 297 2447 300
rect 2416 252 2420 297
rect 2443 244 2447 297
rect 2773 272 2892 275
rect 2777 248 2782 272
rect 2849 250 2853 272
rect 2365 239 2386 243
rect 2377 215 2383 239
rect 2886 248 2892 272
rect 3013 274 3016 280
rect 3013 271 3050 274
rect 3047 268 3050 271
rect 3047 265 3068 268
rect 3077 252 3080 262
rect 3212 259 3216 304
rect 3014 249 3080 252
rect 3239 251 3243 304
rect 2883 244 2904 248
rect 2416 215 2420 237
rect 2487 215 2492 239
rect 2377 212 2496 215
rect 2822 190 2826 243
rect 2849 190 2853 235
rect 3014 231 3017 249
rect 3161 246 3182 250
rect 3173 222 3179 246
rect 3212 222 3216 244
rect 3283 222 3288 246
rect 3173 219 3292 222
rect 2822 187 2853 190
rect 3217 157 3248 160
rect 3018 125 3021 131
rect 3018 122 3055 125
rect 3052 119 3055 122
rect 3052 116 3073 119
rect 3082 103 3085 113
rect 3217 112 3221 157
rect 3244 104 3248 157
rect 3019 100 3085 103
rect 3019 82 3022 100
rect 3166 99 3187 103
rect 3178 75 3184 99
rect 3217 75 3221 97
rect 3288 75 3293 99
rect 3178 72 3297 75
<< m3contact >>
rect 2340 632 2345 637
rect 3159 618 3164 623
rect 2634 550 2639 555
rect 2558 545 2563 550
rect 2780 539 2785 544
rect 2814 540 2819 545
rect 2835 540 2840 545
rect 2857 540 2862 545
rect 2885 541 2890 546
rect 2904 538 2909 544
rect 2337 531 2342 536
rect 2634 476 2639 481
rect 2558 471 2563 476
rect 2336 434 2341 439
rect 2634 407 2639 412
rect 2558 402 2563 407
rect 2337 338 2342 343
rect 2634 333 2639 338
rect 2920 334 2925 339
rect 2558 328 2563 333
<< m123contact >>
rect 2778 725 2783 730
rect 2913 725 2918 730
rect 3051 724 3056 729
rect 2638 708 2643 713
rect 2778 672 2783 677
rect 2796 676 2801 681
rect 2913 672 2918 677
rect 2931 676 2936 681
rect 3051 671 3056 676
rect 3069 675 3074 680
rect 2638 655 2643 660
rect 2656 659 2661 664
rect 2810 631 2815 636
rect 2945 631 2950 636
rect 3083 630 3088 635
rect 2670 614 2675 619
rect 3000 581 3005 586
rect 3000 528 3005 533
rect 3018 532 3023 537
rect 3032 487 3037 492
rect 3011 445 3016 450
rect 3011 392 3016 397
rect 3029 396 3034 401
rect 3043 351 3048 356
rect 3020 311 3025 316
rect 3020 258 3025 263
rect 3038 262 3043 267
rect 3052 217 3057 222
rect 3025 162 3030 167
rect 3025 109 3030 114
rect 3043 113 3048 118
rect 3057 68 3062 73
<< metal3 >>
rect 2638 660 2641 708
rect 2778 677 2781 725
rect 2801 676 2813 679
rect 2661 659 2673 662
rect 2345 632 2356 637
rect 2351 603 2356 632
rect 2670 619 2673 659
rect 2810 636 2813 676
rect 2913 677 2916 725
rect 2936 676 2948 679
rect 2945 636 2948 676
rect 3051 676 3054 724
rect 3074 675 3086 678
rect 3083 635 3086 675
rect 3096 618 3159 623
rect 3096 614 3101 618
rect 3032 609 3101 614
rect 3032 605 3037 609
rect 2351 598 2551 603
rect 2546 550 2551 598
rect 2752 600 3037 605
rect 2752 562 2757 600
rect 2752 557 2769 562
rect 2639 550 2656 555
rect 2546 545 2558 550
rect 2342 531 2353 536
rect 2347 506 2352 531
rect 2651 519 2656 550
rect 2764 554 2769 557
rect 2764 549 2778 554
rect 2773 544 2778 549
rect 2773 539 2780 544
rect 2808 540 2814 545
rect 2808 519 2813 540
rect 2835 535 2839 540
rect 2651 514 2813 519
rect 2347 501 2556 506
rect 2551 476 2556 501
rect 2834 481 2839 535
rect 2639 476 2839 481
rect 2551 471 2558 476
rect 2341 434 2352 439
rect 2347 405 2352 434
rect 2857 412 2862 540
rect 2639 407 2862 412
rect 2881 541 2885 546
rect 2542 405 2558 407
rect 2347 402 2558 405
rect 2347 400 2542 402
rect 2342 338 2353 343
rect 2881 338 2886 541
rect 2348 311 2353 338
rect 2639 333 2886 338
rect 2909 339 2914 544
rect 3000 533 3003 581
rect 3023 532 3035 535
rect 3032 492 3035 532
rect 3011 397 3014 445
rect 3034 396 3046 399
rect 3043 356 3046 396
rect 2909 334 2920 339
rect 2909 333 2914 334
rect 2551 328 2558 333
rect 2551 311 2556 328
rect 2348 306 2556 311
rect 3020 263 3023 311
rect 3043 262 3055 265
rect 3052 222 3055 262
rect 3025 114 3028 162
rect 3048 113 3060 116
rect 3057 73 3060 113
<< labels >>
rlabel metal1 2656 608 2660 611 1 gnd
rlabel metal1 2706 614 2709 616 1 gnd
rlabel metal1 2654 664 2655 666 1 gnd
rlabel metal1 2650 708 2653 710 5 vdd
rlabel metal1 2651 654 2654 656 1 vdd
rlabel metal1 2735 643 2739 647 7 p0
rlabel metal1 2627 678 2628 681 1 a0
rlabel metal1 2627 624 2628 627 1 b0
rlabel metal1 2629 553 2630 554 7 g0
rlabel metal1 2566 547 2567 548 3 b0
rlabel metal1 2564 554 2565 555 3 a0
rlabel metal1 2589 521 2589 521 1 gnd!
rlabel metal1 2589 585 2589 585 5 vdd!
rlabel metal1 2629 479 2630 480 7 g1
rlabel metal1 2589 378 2589 378 1 gnd!
rlabel metal1 2589 442 2589 442 5 vdd!
rlabel metal1 2589 304 2589 304 1 gnd!
rlabel metal1 2589 368 2589 368 5 vdd!
rlabel metal1 2564 411 2565 412 3 a2
rlabel metal1 2566 404 2567 405 3 b2
rlabel metal1 2565 337 2566 338 3 a3
rlabel metal1 2566 330 2567 331 3 b3
rlabel metal1 2629 336 2630 337 7 g3
rlabel metal1 2566 473 2567 474 3 b1
rlabel metal1 2565 480 2566 481 3 a1
rlabel metal1 2589 511 2589 511 5 vdd!
rlabel metal1 2589 447 2589 447 1 gnd!
rlabel metal1 2668 540 2669 541 1 cin
rlabel metal1 2689 540 2690 542 1 p0
rlabel metal1 2722 540 2723 541 1 p1
rlabel metal1 2755 540 2756 541 1 p2
rlabel metal1 2786 540 2787 541 1 p3
rlabel metal1 2796 539 2798 541 1 c3b
rlabel metal1 2820 541 2821 542 1 g0
rlabel metal1 2830 540 2832 542 1 c0b
rlabel metal1 2841 541 2842 542 1 g1
rlabel metal1 2851 540 2853 542 1 c1b
rlabel metal1 3018 481 3022 484 1 gnd
rlabel metal1 3068 487 3071 489 1 gnd
rlabel metal1 3016 537 3017 539 1 gnd
rlabel metal1 3012 581 3015 583 5 vdd
rlabel metal1 3013 527 3016 529 1 vdd
rlabel metal1 3029 345 3033 348 1 gnd
rlabel metal1 3079 351 3082 353 1 gnd
rlabel metal1 3027 401 3028 403 1 gnd
rlabel metal1 3023 445 3026 447 5 vdd
rlabel metal1 3024 391 3027 393 1 vdd
rlabel metal1 3038 211 3042 214 1 gnd
rlabel metal1 3088 217 3091 219 1 gnd
rlabel metal1 3036 267 3037 269 1 gnd
rlabel metal1 3032 311 3035 313 5 vdd
rlabel metal1 3033 257 3036 259 1 vdd
rlabel metal1 3043 62 3047 65 1 gnd
rlabel metal1 3093 68 3096 70 1 gnd
rlabel metal1 3041 118 3042 120 1 gnd
rlabel metal1 3037 162 3040 164 5 vdd
rlabel metal1 3038 108 3041 110 1 vdd
rlabel metal1 2989 551 2990 554 1 p0
rlabel metal1 2989 497 2990 500 1 cin
rlabel metal1 3097 516 3101 520 1 s0
rlabel metal1 3000 415 3001 418 1 p1
rlabel metal1 3000 361 3001 364 1 c0
rlabel metal1 3108 380 3112 384 1 s1
rlabel metal1 3009 281 3010 284 1 p2
rlabel metal1 3009 227 3010 230 1 c1
rlabel metal1 3117 246 3121 250 1 s2
rlabel metal1 3014 132 3015 135 1 p3
rlabel metal1 3014 78 3015 81 1 c2
rlabel metal1 3122 97 3126 101 1 s3
rlabel metal1 2629 410 2630 411 7 g2
rlabel metal1 2391 611 2394 612 1 gnd
rlabel metal1 2397 683 2399 684 5 vdd
rlabel metal2 2380 633 2382 634 1 clk
rlabel metal1 2529 635 2532 639 1 a0
rlabel metal1 2378 640 2380 642 1 a0d
rlabel metal1 2393 513 2396 514 1 gnd
rlabel metal1 2399 585 2401 586 5 vdd
rlabel metal2 2382 535 2384 536 1 clk
rlabel metal1 2392 416 2395 417 1 gnd
rlabel metal1 2398 488 2400 489 5 vdd
rlabel metal2 2381 438 2383 439 1 clk
rlabel metal1 2393 320 2396 321 1 gnd
rlabel metal1 2399 392 2401 393 5 vdd
rlabel metal2 2382 342 2384 343 1 clk
rlabel metal1 2196 608 2199 609 1 gnd
rlabel metal1 2202 680 2204 681 5 vdd
rlabel metal2 2185 630 2187 631 1 clk
rlabel metal2 2182 336 2184 337 1 clk
rlabel metal1 2199 386 2201 387 5 vdd
rlabel metal1 2193 314 2196 315 1 gnd
rlabel metal2 2181 432 2183 433 1 clk
rlabel metal1 2198 482 2200 483 5 vdd
rlabel metal1 2192 410 2195 411 1 gnd
rlabel metal2 2182 529 2184 530 1 clk
rlabel metal1 2199 579 2201 580 5 vdd
rlabel metal1 2193 507 2196 508 1 gnd
rlabel metal1 2183 637 2185 639 1 b0d
rlabel metal1 2334 632 2337 636 1 b0
rlabel metal1 2180 536 2182 538 1 b1d
rlabel metal1 2331 531 2334 535 1 b1
rlabel metal1 2179 439 2181 441 1 b2d
rlabel metal1 2330 434 2333 438 1 b2
rlabel metal1 2180 343 2182 345 1 b3d
rlabel metal1 2331 338 2334 342 1 b3
rlabel metal1 2531 537 2534 541 1 a1
rlabel metal1 2380 542 2382 544 1 a1d
rlabel metal1 2379 445 2381 447 1 a2d
rlabel metal1 2530 440 2533 444 1 a2
rlabel metal1 2380 349 2382 351 1 a3d
rlabel metal1 2395 219 2398 220 1 gnd
rlabel metal1 2401 291 2403 292 5 vdd
rlabel metal2 2384 241 2386 242 1 clk
rlabel metal1 2533 243 2536 247 1 cin
rlabel metal1 2382 249 2384 250 1 cind
rlabel metal1 3168 491 3171 492 1 gnd
rlabel metal1 3174 563 3176 564 5 vdd
rlabel metal2 3157 513 3159 514 1 clk
rlabel metal1 3181 349 3184 350 1 gnd
rlabel metal1 3187 421 3189 422 5 vdd
rlabel metal2 3170 371 3172 372 1 clk
rlabel metal1 3191 226 3194 227 1 gnd
rlabel metal1 3197 298 3199 299 5 vdd
rlabel metal2 3180 248 3182 249 1 clk
rlabel metal1 3196 79 3199 80 1 gnd
rlabel metal1 3202 151 3204 152 5 vdd
rlabel metal2 3185 101 3187 102 1 clk
rlabel metal1 3183 108 3185 110 1 s3
rlabel metal1 3334 103 3337 107 7 s3d
rlabel metal1 3329 250 3332 254 1 s2d
rlabel metal1 3178 255 3180 257 1 s2
rlabel metal1 3168 378 3170 380 1 s1
rlabel metal1 3155 520 3158 522 1 s0
rlabel metal1 3305 515 3310 519 1 s0d
rlabel metal1 3319 373 3322 377 1 s1d
rlabel metal1 2844 305 2847 307 1 gnd
rlabel metal1 2775 305 2782 310 1 c2b
rlabel metal1 2740 305 2747 310 1 c1b
rlabel metal1 2701 305 2708 310 1 c0b
rlabel metal1 2673 299 2679 301 1 gnd
rlabel metal1 2531 344 2534 348 1 a3
rlabel metal1 2783 597 2790 598 1 vdd
rlabel metal1 2787 565 2788 566 1 c0b
rlabel metal1 2772 564 2775 566 1 gnd
rlabel metal1 2823 566 2824 567 1 c1b
rlabel metal1 2808 565 2811 567 1 gnd
rlabel metal1 2819 598 2826 599 1 vdd
rlabel metal1 2857 598 2864 599 1 vdd
rlabel metal1 2846 565 2849 567 1 gnd
rlabel metal1 2861 566 2862 567 1 c2b
rlabel metal1 2796 625 2800 628 1 gnd
rlabel metal1 2846 631 2849 633 1 gnd
rlabel metal1 2794 681 2795 683 1 gnd
rlabel metal1 2790 725 2793 727 5 vdd
rlabel metal1 2791 671 2794 673 1 vdd
rlabel metal1 2931 625 2935 628 1 gnd
rlabel metal1 2981 631 2984 633 1 gnd
rlabel metal1 2929 681 2930 683 1 gnd
rlabel metal1 2925 725 2928 727 5 vdd
rlabel metal1 2926 671 2929 673 1 vdd
rlabel metal1 3069 624 3073 627 1 gnd
rlabel metal1 3119 630 3122 632 1 gnd
rlabel metal1 3067 680 3068 682 1 gnd
rlabel metal1 3063 724 3066 726 5 vdd
rlabel metal1 3064 670 3067 672 1 vdd
rlabel metal1 2767 641 2768 644 1 b1
rlabel metal1 2767 695 2768 698 1 a1
rlabel metal1 2902 695 2903 698 1 a2
rlabel metal1 2902 641 2903 644 1 b2
rlabel metal1 3040 694 3041 697 1 a3
rlabel metal1 3040 640 3041 643 1 b3
rlabel metal1 3148 659 3152 663 7 p3
rlabel metal1 2875 660 2879 664 1 p1
rlabel metal1 3010 660 3014 664 1 p2
rlabel metal1 2891 542 2892 543 1 g3
rlabel metal1 2901 541 2903 543 1 c3b
rlabel metal1 2863 541 2864 542 1 g2
rlabel metal1 2873 540 2875 542 1 c2b
rlabel metal1 2937 483 2940 485 1 c1b
rlabel metal1 2960 484 2961 485 1 c1
rlabel metal1 2939 452 2941 453 1 gnd
rlabel metal1 2947 515 2949 516 1 vdd
rlabel metal1 2931 559 2932 561 1 c0b
rlabel metal1 2955 560 2958 562 1 c0
rlabel metal1 2932 528 2934 529 1 gnd
rlabel metal1 2941 591 2943 592 1 vdd
rlabel metal1 2896 597 2903 598 1 vdd
rlabel metal1 2885 564 2888 566 1 gnd
rlabel metal1 2900 565 2901 566 1 c3b
rlabel metal1 2941 407 2944 409 1 c2b
rlabel metal1 2963 408 2964 409 1 c2
rlabel metal1 2942 377 2944 378 1 gnd
rlabel metal1 2948 439 2950 440 1 vdd
rlabel metal1 2930 335 2933 337 1 c3b
rlabel metal1 2952 336 2953 337 1 c3
rlabel metal1 2930 304 2932 305 1 gnd
rlabel metal1 2937 367 2939 368 1 vdd
rlabel metal1 2871 267 2874 268 5 gnd
rlabel metal1 2866 195 2868 196 1 vdd
rlabel metal2 2883 245 2885 246 5 clk
rlabel metal1 2885 237 2887 239 5 c3
rlabel metal1 2733 240 2736 244 5 coutd
<< end >>
