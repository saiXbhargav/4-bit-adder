magic
tech scmos
timestamp 1731695463
<< nwell >>
rect 517 -474 541 -450
rect 556 -460 590 -454
rect 65 -517 97 -480
rect 103 -517 129 -480
rect 147 -517 173 -480
rect 192 -517 218 -480
rect 260 -514 292 -477
rect 298 -514 324 -477
rect 342 -514 368 -477
rect 387 -514 413 -477
rect 556 -490 618 -460
rect 657 -474 681 -450
rect 696 -460 730 -454
rect 696 -490 758 -460
rect 792 -474 816 -450
rect 831 -460 865 -454
rect 831 -490 893 -460
rect 930 -475 954 -451
rect 969 -461 1003 -455
rect 584 -496 618 -490
rect 724 -496 758 -490
rect 859 -496 893 -490
rect 969 -491 1031 -461
rect 997 -497 1031 -491
rect 517 -529 541 -505
rect 657 -529 681 -505
rect 792 -529 816 -505
rect 930 -530 954 -506
rect 62 -618 94 -581
rect 100 -618 126 -581
rect 144 -618 170 -581
rect 189 -618 215 -581
rect 262 -612 294 -575
rect 300 -612 326 -575
rect 344 -612 370 -575
rect 389 -612 415 -575
rect 442 -601 479 -575
rect 485 -601 513 -575
rect 548 -599 576 -573
rect 584 -599 612 -573
rect 625 -599 653 -573
rect 660 -599 688 -573
rect 794 -624 822 -598
rect 879 -601 903 -577
rect 918 -587 952 -581
rect 918 -617 980 -587
rect 946 -623 980 -617
rect 61 -715 93 -678
rect 99 -715 125 -678
rect 143 -715 169 -678
rect 188 -715 214 -678
rect 261 -709 293 -672
rect 299 -709 325 -672
rect 343 -709 369 -672
rect 388 -709 414 -672
rect 442 -675 479 -649
rect 485 -675 513 -649
rect 879 -656 903 -632
rect 1037 -634 1069 -597
rect 1075 -634 1101 -597
rect 1119 -634 1145 -597
rect 1164 -634 1190 -597
rect 795 -709 823 -683
rect 442 -744 479 -718
rect 485 -744 513 -718
rect 890 -737 914 -713
rect 929 -723 963 -717
rect 929 -753 991 -723
rect 957 -759 991 -753
rect 62 -811 94 -774
rect 100 -811 126 -774
rect 144 -811 170 -774
rect 189 -811 215 -774
rect 262 -805 294 -768
rect 300 -805 326 -768
rect 344 -805 370 -768
rect 389 -805 415 -768
rect 890 -792 914 -768
rect 1050 -776 1082 -739
rect 1088 -776 1114 -739
rect 1132 -776 1158 -739
rect 1177 -776 1203 -739
rect 442 -818 479 -792
rect 485 -818 513 -792
rect 798 -820 826 -794
rect 264 -906 296 -869
rect 302 -906 328 -869
rect 346 -906 372 -869
rect 391 -906 417 -869
rect 799 -892 827 -866
rect 899 -871 923 -847
rect 938 -857 972 -851
rect 938 -887 1000 -857
rect 966 -893 1000 -887
rect 1060 -899 1092 -862
rect 1098 -899 1124 -862
rect 1142 -899 1168 -862
rect 1187 -899 1213 -862
rect 899 -926 923 -902
rect 629 -975 661 -938
rect 667 -975 693 -938
rect 711 -975 737 -938
rect 756 -975 782 -938
rect 904 -1020 928 -996
rect 943 -1006 977 -1000
rect 943 -1036 1005 -1006
rect 971 -1042 1005 -1036
rect 1065 -1046 1097 -1009
rect 1103 -1046 1129 -1009
rect 1147 -1046 1173 -1009
rect 1192 -1046 1218 -1009
rect 904 -1075 928 -1051
<< ntransistor >>
rect 528 -488 530 -482
rect 668 -488 670 -482
rect 72 -543 74 -533
rect 108 -543 110 -533
rect 116 -543 118 -533
rect 152 -543 154 -533
rect 160 -543 162 -533
rect 203 -543 205 -533
rect 267 -540 269 -530
rect 303 -540 305 -530
rect 311 -540 313 -530
rect 347 -540 349 -530
rect 355 -540 357 -530
rect 398 -540 400 -530
rect 803 -488 805 -482
rect 567 -537 569 -525
rect 577 -537 579 -525
rect 595 -537 597 -525
rect 605 -537 607 -525
rect 941 -489 943 -483
rect 707 -537 709 -525
rect 717 -537 719 -525
rect 735 -537 737 -525
rect 745 -537 747 -525
rect 842 -537 844 -525
rect 852 -537 854 -525
rect 870 -537 872 -525
rect 880 -537 882 -525
rect 528 -543 530 -537
rect 668 -543 670 -537
rect 803 -543 805 -537
rect 980 -538 982 -526
rect 990 -538 992 -526
rect 1008 -538 1010 -526
rect 1018 -538 1020 -526
rect 941 -544 943 -538
rect 69 -644 71 -634
rect 105 -644 107 -634
rect 113 -644 115 -634
rect 149 -644 151 -634
rect 157 -644 159 -634
rect 200 -644 202 -634
rect 269 -638 271 -628
rect 305 -638 307 -628
rect 313 -638 315 -628
rect 349 -638 351 -628
rect 357 -638 359 -628
rect 400 -638 402 -628
rect 455 -629 457 -616
rect 465 -629 467 -616
rect 497 -618 499 -611
rect 890 -615 892 -609
rect 455 -703 457 -690
rect 465 -703 467 -690
rect 497 -692 499 -685
rect 68 -741 70 -731
rect 104 -741 106 -731
rect 112 -741 114 -731
rect 148 -741 150 -731
rect 156 -741 158 -731
rect 199 -741 201 -731
rect 268 -735 270 -725
rect 304 -735 306 -725
rect 312 -735 314 -725
rect 348 -735 350 -725
rect 356 -735 358 -725
rect 399 -735 401 -725
rect 455 -772 457 -759
rect 465 -772 467 -759
rect 497 -761 499 -754
rect 69 -837 71 -827
rect 105 -837 107 -827
rect 113 -837 115 -827
rect 149 -837 151 -827
rect 157 -837 159 -827
rect 200 -837 202 -827
rect 269 -831 271 -821
rect 305 -831 307 -821
rect 313 -831 315 -821
rect 349 -831 351 -821
rect 357 -831 359 -821
rect 400 -831 402 -821
rect 455 -846 457 -833
rect 465 -846 467 -833
rect 497 -835 499 -828
rect 553 -847 555 -623
rect 560 -847 562 -623
rect 607 -846 609 -622
rect 640 -846 642 -622
rect 671 -846 673 -622
rect 705 -845 707 -621
rect 726 -845 728 -621
rect 743 -845 745 -621
rect 761 -844 763 -620
rect 806 -641 808 -634
rect 929 -664 931 -652
rect 939 -664 941 -652
rect 957 -664 959 -652
rect 967 -664 969 -652
rect 1044 -660 1046 -650
rect 1080 -660 1082 -650
rect 1088 -660 1090 -650
rect 1124 -660 1126 -650
rect 1132 -660 1134 -650
rect 1175 -660 1177 -650
rect 890 -670 892 -664
rect 807 -726 809 -719
rect 901 -751 903 -745
rect 940 -800 942 -788
rect 950 -800 952 -788
rect 968 -800 970 -788
rect 978 -800 980 -788
rect 901 -806 903 -800
rect 1057 -802 1059 -792
rect 1093 -802 1095 -792
rect 1101 -802 1103 -792
rect 1137 -802 1139 -792
rect 1145 -802 1147 -792
rect 1188 -802 1190 -792
rect 810 -837 812 -830
rect 910 -885 912 -879
rect 811 -909 813 -902
rect 271 -932 273 -922
rect 307 -932 309 -922
rect 315 -932 317 -922
rect 351 -932 353 -922
rect 359 -932 361 -922
rect 402 -932 404 -922
rect 949 -934 951 -922
rect 959 -934 961 -922
rect 977 -934 979 -922
rect 987 -934 989 -922
rect 1067 -925 1069 -915
rect 1103 -925 1105 -915
rect 1111 -925 1113 -915
rect 1147 -925 1149 -915
rect 1155 -925 1157 -915
rect 1198 -925 1200 -915
rect 910 -940 912 -934
rect 636 -1001 638 -991
rect 672 -1001 674 -991
rect 680 -1001 682 -991
rect 716 -1001 718 -991
rect 724 -1001 726 -991
rect 767 -1001 769 -991
rect 915 -1034 917 -1028
rect 954 -1083 956 -1071
rect 964 -1083 966 -1071
rect 982 -1083 984 -1071
rect 992 -1083 994 -1071
rect 1072 -1072 1074 -1062
rect 1108 -1072 1110 -1062
rect 1116 -1072 1118 -1062
rect 1152 -1072 1154 -1062
rect 1160 -1072 1162 -1062
rect 1203 -1072 1205 -1062
rect 915 -1089 917 -1083
<< ptransistor >>
rect 528 -468 530 -456
rect 76 -511 78 -486
rect 84 -511 86 -486
rect 114 -511 116 -486
rect 158 -511 160 -486
rect 203 -511 205 -486
rect 271 -508 273 -483
rect 279 -508 281 -483
rect 309 -508 311 -483
rect 353 -508 355 -483
rect 398 -508 400 -483
rect 567 -484 569 -460
rect 577 -484 579 -460
rect 595 -490 597 -466
rect 605 -490 607 -466
rect 668 -468 670 -456
rect 707 -484 709 -460
rect 717 -484 719 -460
rect 528 -523 530 -511
rect 735 -490 737 -466
rect 745 -490 747 -466
rect 803 -468 805 -456
rect 842 -484 844 -460
rect 852 -484 854 -460
rect 668 -523 670 -511
rect 870 -490 872 -466
rect 880 -490 882 -466
rect 941 -469 943 -457
rect 980 -485 982 -461
rect 990 -485 992 -461
rect 803 -523 805 -511
rect 1008 -491 1010 -467
rect 1018 -491 1020 -467
rect 941 -524 943 -512
rect 73 -612 75 -587
rect 81 -612 83 -587
rect 111 -612 113 -587
rect 155 -612 157 -587
rect 200 -612 202 -587
rect 273 -606 275 -581
rect 281 -606 283 -581
rect 311 -606 313 -581
rect 355 -606 357 -581
rect 400 -606 402 -581
rect 455 -593 457 -581
rect 465 -593 467 -581
rect 497 -593 499 -581
rect 560 -591 562 -579
rect 596 -591 598 -579
rect 637 -591 639 -579
rect 672 -591 674 -579
rect 890 -595 892 -583
rect 806 -616 808 -604
rect 929 -611 931 -587
rect 939 -611 941 -587
rect 455 -667 457 -655
rect 465 -667 467 -655
rect 497 -667 499 -655
rect 72 -709 74 -684
rect 80 -709 82 -684
rect 110 -709 112 -684
rect 154 -709 156 -684
rect 199 -709 201 -684
rect 272 -703 274 -678
rect 280 -703 282 -678
rect 310 -703 312 -678
rect 354 -703 356 -678
rect 399 -703 401 -678
rect 455 -736 457 -724
rect 465 -736 467 -724
rect 497 -736 499 -724
rect 73 -805 75 -780
rect 81 -805 83 -780
rect 111 -805 113 -780
rect 155 -805 157 -780
rect 200 -805 202 -780
rect 273 -799 275 -774
rect 281 -799 283 -774
rect 311 -799 313 -774
rect 355 -799 357 -774
rect 400 -799 402 -774
rect 455 -810 457 -798
rect 465 -810 467 -798
rect 497 -810 499 -798
rect 957 -617 959 -593
rect 967 -617 969 -593
rect 890 -650 892 -638
rect 1048 -628 1050 -603
rect 1056 -628 1058 -603
rect 1086 -628 1088 -603
rect 1130 -628 1132 -603
rect 1175 -628 1177 -603
rect 807 -701 809 -689
rect 901 -731 903 -719
rect 940 -747 942 -723
rect 950 -747 952 -723
rect 968 -753 970 -729
rect 978 -753 980 -729
rect 901 -786 903 -774
rect 1061 -770 1063 -745
rect 1069 -770 1071 -745
rect 1099 -770 1101 -745
rect 1143 -770 1145 -745
rect 1188 -770 1190 -745
rect 810 -812 812 -800
rect 910 -865 912 -853
rect 275 -900 277 -875
rect 283 -900 285 -875
rect 313 -900 315 -875
rect 357 -900 359 -875
rect 402 -900 404 -875
rect 811 -884 813 -872
rect 949 -881 951 -857
rect 959 -881 961 -857
rect 977 -887 979 -863
rect 987 -887 989 -863
rect 910 -920 912 -908
rect 1071 -893 1073 -868
rect 1079 -893 1081 -868
rect 1109 -893 1111 -868
rect 1153 -893 1155 -868
rect 1198 -893 1200 -868
rect 640 -969 642 -944
rect 648 -969 650 -944
rect 678 -969 680 -944
rect 722 -969 724 -944
rect 767 -969 769 -944
rect 915 -1014 917 -1002
rect 954 -1030 956 -1006
rect 964 -1030 966 -1006
rect 982 -1036 984 -1012
rect 992 -1036 994 -1012
rect 915 -1069 917 -1057
rect 1076 -1040 1078 -1015
rect 1084 -1040 1086 -1015
rect 1114 -1040 1116 -1015
rect 1158 -1040 1160 -1015
rect 1203 -1040 1205 -1015
<< ndiffusion >>
rect 527 -488 528 -482
rect 530 -488 531 -482
rect 667 -488 668 -482
rect 670 -488 671 -482
rect 71 -543 72 -533
rect 74 -543 75 -533
rect 107 -543 108 -533
rect 110 -543 111 -533
rect 115 -543 116 -533
rect 118 -543 119 -533
rect 151 -543 152 -533
rect 154 -543 155 -533
rect 159 -543 160 -533
rect 162 -543 163 -533
rect 202 -543 203 -533
rect 205 -543 206 -533
rect 266 -540 267 -530
rect 269 -540 270 -530
rect 302 -540 303 -530
rect 305 -540 306 -530
rect 310 -540 311 -530
rect 313 -540 314 -530
rect 346 -540 347 -530
rect 349 -540 350 -530
rect 354 -540 355 -530
rect 357 -540 358 -530
rect 397 -540 398 -530
rect 400 -540 401 -530
rect 802 -488 803 -482
rect 805 -488 806 -482
rect 566 -537 567 -525
rect 569 -537 577 -525
rect 579 -537 580 -525
rect 594 -537 595 -525
rect 597 -537 605 -525
rect 607 -537 608 -525
rect 940 -489 941 -483
rect 943 -489 944 -483
rect 706 -537 707 -525
rect 709 -537 717 -525
rect 719 -537 720 -525
rect 734 -537 735 -525
rect 737 -537 745 -525
rect 747 -537 748 -525
rect 841 -537 842 -525
rect 844 -537 852 -525
rect 854 -537 855 -525
rect 869 -537 870 -525
rect 872 -537 880 -525
rect 882 -537 883 -525
rect 527 -543 528 -537
rect 530 -543 531 -537
rect 667 -543 668 -537
rect 670 -543 671 -537
rect 802 -543 803 -537
rect 805 -543 806 -537
rect 979 -538 980 -526
rect 982 -538 990 -526
rect 992 -538 993 -526
rect 1007 -538 1008 -526
rect 1010 -538 1018 -526
rect 1020 -538 1021 -526
rect 940 -544 941 -538
rect 943 -544 944 -538
rect 68 -644 69 -634
rect 71 -644 72 -634
rect 104 -644 105 -634
rect 107 -644 108 -634
rect 112 -644 113 -634
rect 115 -644 116 -634
rect 148 -644 149 -634
rect 151 -644 152 -634
rect 156 -644 157 -634
rect 159 -644 160 -634
rect 199 -644 200 -634
rect 202 -644 203 -634
rect 268 -638 269 -628
rect 271 -638 272 -628
rect 304 -638 305 -628
rect 307 -638 308 -628
rect 312 -638 313 -628
rect 315 -638 316 -628
rect 348 -638 349 -628
rect 351 -638 352 -628
rect 356 -638 357 -628
rect 359 -638 360 -628
rect 399 -638 400 -628
rect 402 -638 403 -628
rect 454 -629 455 -616
rect 457 -629 465 -616
rect 467 -629 468 -616
rect 496 -618 497 -611
rect 499 -618 500 -611
rect 889 -615 890 -609
rect 892 -615 893 -609
rect 454 -703 455 -690
rect 457 -703 465 -690
rect 467 -703 468 -690
rect 496 -692 497 -685
rect 499 -692 500 -685
rect 67 -741 68 -731
rect 70 -741 71 -731
rect 103 -741 104 -731
rect 106 -741 107 -731
rect 111 -741 112 -731
rect 114 -741 115 -731
rect 147 -741 148 -731
rect 150 -741 151 -731
rect 155 -741 156 -731
rect 158 -741 159 -731
rect 198 -741 199 -731
rect 201 -741 202 -731
rect 267 -735 268 -725
rect 270 -735 271 -725
rect 303 -735 304 -725
rect 306 -735 307 -725
rect 311 -735 312 -725
rect 314 -735 315 -725
rect 347 -735 348 -725
rect 350 -735 351 -725
rect 355 -735 356 -725
rect 358 -735 359 -725
rect 398 -735 399 -725
rect 401 -735 402 -725
rect 454 -772 455 -759
rect 457 -772 465 -759
rect 467 -772 468 -759
rect 496 -761 497 -754
rect 499 -761 500 -754
rect 68 -837 69 -827
rect 71 -837 72 -827
rect 104 -837 105 -827
rect 107 -837 108 -827
rect 112 -837 113 -827
rect 115 -837 116 -827
rect 148 -837 149 -827
rect 151 -837 152 -827
rect 156 -837 157 -827
rect 159 -837 160 -827
rect 199 -837 200 -827
rect 202 -837 203 -827
rect 268 -831 269 -821
rect 271 -831 272 -821
rect 304 -831 305 -821
rect 307 -831 308 -821
rect 312 -831 313 -821
rect 315 -831 316 -821
rect 348 -831 349 -821
rect 351 -831 352 -821
rect 356 -831 357 -821
rect 359 -831 360 -821
rect 399 -831 400 -821
rect 402 -831 403 -821
rect 454 -846 455 -833
rect 457 -846 465 -833
rect 467 -846 468 -833
rect 496 -835 497 -828
rect 499 -835 500 -828
rect 552 -847 553 -623
rect 555 -847 560 -623
rect 562 -847 563 -623
rect 606 -846 607 -622
rect 609 -846 610 -622
rect 639 -846 640 -622
rect 642 -846 643 -622
rect 670 -846 671 -622
rect 673 -846 674 -622
rect 704 -845 705 -621
rect 707 -845 708 -621
rect 725 -845 726 -621
rect 728 -845 729 -621
rect 742 -845 743 -621
rect 745 -845 746 -621
rect 760 -844 761 -620
rect 763 -844 764 -620
rect 805 -641 806 -634
rect 808 -641 809 -634
rect 928 -664 929 -652
rect 931 -664 939 -652
rect 941 -664 942 -652
rect 956 -664 957 -652
rect 959 -664 967 -652
rect 969 -664 970 -652
rect 1043 -660 1044 -650
rect 1046 -660 1047 -650
rect 1079 -660 1080 -650
rect 1082 -660 1083 -650
rect 1087 -660 1088 -650
rect 1090 -660 1091 -650
rect 1123 -660 1124 -650
rect 1126 -660 1127 -650
rect 1131 -660 1132 -650
rect 1134 -660 1135 -650
rect 1174 -660 1175 -650
rect 1177 -660 1178 -650
rect 889 -670 890 -664
rect 892 -670 893 -664
rect 806 -726 807 -719
rect 809 -726 810 -719
rect 900 -751 901 -745
rect 903 -751 904 -745
rect 939 -800 940 -788
rect 942 -800 950 -788
rect 952 -800 953 -788
rect 967 -800 968 -788
rect 970 -800 978 -788
rect 980 -800 981 -788
rect 900 -806 901 -800
rect 903 -806 904 -800
rect 1056 -802 1057 -792
rect 1059 -802 1060 -792
rect 1092 -802 1093 -792
rect 1095 -802 1096 -792
rect 1100 -802 1101 -792
rect 1103 -802 1104 -792
rect 1136 -802 1137 -792
rect 1139 -802 1140 -792
rect 1144 -802 1145 -792
rect 1147 -802 1148 -792
rect 1187 -802 1188 -792
rect 1190 -802 1191 -792
rect 809 -837 810 -830
rect 812 -837 813 -830
rect 909 -885 910 -879
rect 912 -885 913 -879
rect 810 -909 811 -902
rect 813 -909 814 -902
rect 270 -932 271 -922
rect 273 -932 274 -922
rect 306 -932 307 -922
rect 309 -932 310 -922
rect 314 -932 315 -922
rect 317 -932 318 -922
rect 350 -932 351 -922
rect 353 -932 354 -922
rect 358 -932 359 -922
rect 361 -932 362 -922
rect 401 -932 402 -922
rect 404 -932 405 -922
rect 948 -934 949 -922
rect 951 -934 959 -922
rect 961 -934 962 -922
rect 976 -934 977 -922
rect 979 -934 987 -922
rect 989 -934 990 -922
rect 1066 -925 1067 -915
rect 1069 -925 1070 -915
rect 1102 -925 1103 -915
rect 1105 -925 1106 -915
rect 1110 -925 1111 -915
rect 1113 -925 1114 -915
rect 1146 -925 1147 -915
rect 1149 -925 1150 -915
rect 1154 -925 1155 -915
rect 1157 -925 1158 -915
rect 1197 -925 1198 -915
rect 1200 -925 1201 -915
rect 909 -940 910 -934
rect 912 -940 913 -934
rect 635 -1001 636 -991
rect 638 -1001 639 -991
rect 671 -1001 672 -991
rect 674 -1001 675 -991
rect 679 -1001 680 -991
rect 682 -1001 683 -991
rect 715 -1001 716 -991
rect 718 -1001 719 -991
rect 723 -1001 724 -991
rect 726 -1001 727 -991
rect 766 -1001 767 -991
rect 769 -1001 770 -991
rect 914 -1034 915 -1028
rect 917 -1034 918 -1028
rect 953 -1083 954 -1071
rect 956 -1083 964 -1071
rect 966 -1083 967 -1071
rect 981 -1083 982 -1071
rect 984 -1083 992 -1071
rect 994 -1083 995 -1071
rect 1071 -1072 1072 -1062
rect 1074 -1072 1075 -1062
rect 1107 -1072 1108 -1062
rect 1110 -1072 1111 -1062
rect 1115 -1072 1116 -1062
rect 1118 -1072 1119 -1062
rect 1151 -1072 1152 -1062
rect 1154 -1072 1155 -1062
rect 1159 -1072 1160 -1062
rect 1162 -1072 1163 -1062
rect 1202 -1072 1203 -1062
rect 1205 -1072 1206 -1062
rect 914 -1089 915 -1083
rect 917 -1089 918 -1083
<< pdiffusion >>
rect 527 -468 528 -456
rect 530 -468 531 -456
rect 75 -511 76 -486
rect 78 -511 79 -486
rect 83 -511 84 -486
rect 86 -511 87 -486
rect 113 -511 114 -486
rect 116 -511 117 -486
rect 157 -511 158 -486
rect 160 -511 161 -486
rect 202 -511 203 -486
rect 205 -511 206 -486
rect 270 -508 271 -483
rect 273 -508 274 -483
rect 278 -508 279 -483
rect 281 -508 282 -483
rect 308 -508 309 -483
rect 311 -508 312 -483
rect 352 -508 353 -483
rect 355 -508 356 -483
rect 397 -508 398 -483
rect 400 -508 401 -483
rect 566 -484 567 -460
rect 569 -484 571 -460
rect 575 -484 577 -460
rect 579 -484 580 -460
rect 594 -490 595 -466
rect 597 -490 599 -466
rect 603 -490 605 -466
rect 607 -490 608 -466
rect 667 -468 668 -456
rect 670 -468 671 -456
rect 706 -484 707 -460
rect 709 -484 711 -460
rect 715 -484 717 -460
rect 719 -484 720 -460
rect 527 -523 528 -511
rect 530 -523 531 -511
rect 734 -490 735 -466
rect 737 -490 739 -466
rect 743 -490 745 -466
rect 747 -490 748 -466
rect 802 -468 803 -456
rect 805 -468 806 -456
rect 841 -484 842 -460
rect 844 -484 846 -460
rect 850 -484 852 -460
rect 854 -484 855 -460
rect 667 -523 668 -511
rect 670 -523 671 -511
rect 869 -490 870 -466
rect 872 -490 874 -466
rect 878 -490 880 -466
rect 882 -490 883 -466
rect 940 -469 941 -457
rect 943 -469 944 -457
rect 979 -485 980 -461
rect 982 -485 984 -461
rect 988 -485 990 -461
rect 992 -485 993 -461
rect 802 -523 803 -511
rect 805 -523 806 -511
rect 1007 -491 1008 -467
rect 1010 -491 1012 -467
rect 1016 -491 1018 -467
rect 1020 -491 1021 -467
rect 940 -524 941 -512
rect 943 -524 944 -512
rect 72 -612 73 -587
rect 75 -612 76 -587
rect 80 -612 81 -587
rect 83 -612 84 -587
rect 110 -612 111 -587
rect 113 -612 114 -587
rect 154 -612 155 -587
rect 157 -612 158 -587
rect 199 -612 200 -587
rect 202 -612 203 -587
rect 272 -606 273 -581
rect 275 -606 276 -581
rect 280 -606 281 -581
rect 283 -606 284 -581
rect 310 -606 311 -581
rect 313 -606 314 -581
rect 354 -606 355 -581
rect 357 -606 358 -581
rect 399 -606 400 -581
rect 402 -606 403 -581
rect 454 -593 455 -581
rect 457 -593 459 -581
rect 463 -593 465 -581
rect 467 -593 468 -581
rect 496 -593 497 -581
rect 499 -593 500 -581
rect 559 -591 560 -579
rect 562 -591 563 -579
rect 595 -591 596 -579
rect 598 -591 599 -579
rect 636 -591 637 -579
rect 639 -591 640 -579
rect 671 -591 672 -579
rect 674 -591 675 -579
rect 889 -595 890 -583
rect 892 -595 893 -583
rect 805 -616 806 -604
rect 808 -616 809 -604
rect 928 -611 929 -587
rect 931 -611 933 -587
rect 937 -611 939 -587
rect 941 -611 942 -587
rect 454 -667 455 -655
rect 457 -667 459 -655
rect 463 -667 465 -655
rect 467 -667 468 -655
rect 496 -667 497 -655
rect 499 -667 500 -655
rect 71 -709 72 -684
rect 74 -709 75 -684
rect 79 -709 80 -684
rect 82 -709 83 -684
rect 109 -709 110 -684
rect 112 -709 113 -684
rect 153 -709 154 -684
rect 156 -709 157 -684
rect 198 -709 199 -684
rect 201 -709 202 -684
rect 271 -703 272 -678
rect 274 -703 275 -678
rect 279 -703 280 -678
rect 282 -703 283 -678
rect 309 -703 310 -678
rect 312 -703 313 -678
rect 353 -703 354 -678
rect 356 -703 357 -678
rect 398 -703 399 -678
rect 401 -703 402 -678
rect 454 -736 455 -724
rect 457 -736 459 -724
rect 463 -736 465 -724
rect 467 -736 468 -724
rect 496 -736 497 -724
rect 499 -736 500 -724
rect 72 -805 73 -780
rect 75 -805 76 -780
rect 80 -805 81 -780
rect 83 -805 84 -780
rect 110 -805 111 -780
rect 113 -805 114 -780
rect 154 -805 155 -780
rect 157 -805 158 -780
rect 199 -805 200 -780
rect 202 -805 203 -780
rect 272 -799 273 -774
rect 275 -799 276 -774
rect 280 -799 281 -774
rect 283 -799 284 -774
rect 310 -799 311 -774
rect 313 -799 314 -774
rect 354 -799 355 -774
rect 357 -799 358 -774
rect 399 -799 400 -774
rect 402 -799 403 -774
rect 454 -810 455 -798
rect 457 -810 459 -798
rect 463 -810 465 -798
rect 467 -810 468 -798
rect 496 -810 497 -798
rect 499 -810 500 -798
rect 956 -617 957 -593
rect 959 -617 961 -593
rect 965 -617 967 -593
rect 969 -617 970 -593
rect 889 -650 890 -638
rect 892 -650 893 -638
rect 1047 -628 1048 -603
rect 1050 -628 1051 -603
rect 1055 -628 1056 -603
rect 1058 -628 1059 -603
rect 1085 -628 1086 -603
rect 1088 -628 1089 -603
rect 1129 -628 1130 -603
rect 1132 -628 1133 -603
rect 1174 -628 1175 -603
rect 1177 -628 1178 -603
rect 806 -701 807 -689
rect 809 -701 810 -689
rect 900 -731 901 -719
rect 903 -731 904 -719
rect 939 -747 940 -723
rect 942 -747 944 -723
rect 948 -747 950 -723
rect 952 -747 953 -723
rect 967 -753 968 -729
rect 970 -753 972 -729
rect 976 -753 978 -729
rect 980 -753 981 -729
rect 900 -786 901 -774
rect 903 -786 904 -774
rect 1060 -770 1061 -745
rect 1063 -770 1064 -745
rect 1068 -770 1069 -745
rect 1071 -770 1072 -745
rect 1098 -770 1099 -745
rect 1101 -770 1102 -745
rect 1142 -770 1143 -745
rect 1145 -770 1146 -745
rect 1187 -770 1188 -745
rect 1190 -770 1191 -745
rect 809 -812 810 -800
rect 812 -812 813 -800
rect 909 -865 910 -853
rect 912 -865 913 -853
rect 274 -900 275 -875
rect 277 -900 278 -875
rect 282 -900 283 -875
rect 285 -900 286 -875
rect 312 -900 313 -875
rect 315 -900 316 -875
rect 356 -900 357 -875
rect 359 -900 360 -875
rect 401 -900 402 -875
rect 404 -900 405 -875
rect 810 -884 811 -872
rect 813 -884 814 -872
rect 948 -881 949 -857
rect 951 -881 953 -857
rect 957 -881 959 -857
rect 961 -881 962 -857
rect 976 -887 977 -863
rect 979 -887 981 -863
rect 985 -887 987 -863
rect 989 -887 990 -863
rect 909 -920 910 -908
rect 912 -920 913 -908
rect 1070 -893 1071 -868
rect 1073 -893 1074 -868
rect 1078 -893 1079 -868
rect 1081 -893 1082 -868
rect 1108 -893 1109 -868
rect 1111 -893 1112 -868
rect 1152 -893 1153 -868
rect 1155 -893 1156 -868
rect 1197 -893 1198 -868
rect 1200 -893 1201 -868
rect 639 -969 640 -944
rect 642 -969 643 -944
rect 647 -969 648 -944
rect 650 -969 651 -944
rect 677 -969 678 -944
rect 680 -969 681 -944
rect 721 -969 722 -944
rect 724 -969 725 -944
rect 766 -969 767 -944
rect 769 -969 770 -944
rect 914 -1014 915 -1002
rect 917 -1014 918 -1002
rect 953 -1030 954 -1006
rect 956 -1030 958 -1006
rect 962 -1030 964 -1006
rect 966 -1030 967 -1006
rect 981 -1036 982 -1012
rect 984 -1036 986 -1012
rect 990 -1036 992 -1012
rect 994 -1036 995 -1012
rect 914 -1069 915 -1057
rect 917 -1069 918 -1057
rect 1075 -1040 1076 -1015
rect 1078 -1040 1079 -1015
rect 1083 -1040 1084 -1015
rect 1086 -1040 1087 -1015
rect 1113 -1040 1114 -1015
rect 1116 -1040 1117 -1015
rect 1157 -1040 1158 -1015
rect 1160 -1040 1161 -1015
rect 1202 -1040 1203 -1015
rect 1205 -1040 1206 -1015
<< ndcontact >>
rect 523 -488 527 -482
rect 531 -488 535 -482
rect 663 -488 667 -482
rect 671 -488 675 -482
rect 67 -543 71 -533
rect 75 -543 79 -533
rect 103 -543 107 -533
rect 111 -543 115 -533
rect 119 -543 123 -533
rect 147 -543 151 -533
rect 155 -543 159 -533
rect 163 -543 167 -533
rect 198 -543 202 -533
rect 206 -543 210 -533
rect 262 -540 266 -530
rect 270 -540 274 -530
rect 298 -540 302 -530
rect 306 -540 310 -530
rect 314 -540 318 -530
rect 342 -540 346 -530
rect 350 -540 354 -530
rect 358 -540 362 -530
rect 393 -540 397 -530
rect 401 -540 405 -530
rect 798 -488 802 -482
rect 806 -488 810 -482
rect 562 -537 566 -525
rect 580 -537 584 -525
rect 590 -537 594 -525
rect 608 -537 612 -525
rect 936 -489 940 -483
rect 944 -489 948 -483
rect 702 -537 706 -525
rect 720 -537 724 -525
rect 730 -537 734 -525
rect 748 -537 752 -525
rect 837 -537 841 -525
rect 855 -537 859 -525
rect 865 -537 869 -525
rect 883 -537 887 -525
rect 523 -543 527 -537
rect 531 -543 535 -537
rect 663 -543 667 -537
rect 671 -543 675 -537
rect 798 -543 802 -537
rect 806 -543 810 -537
rect 975 -538 979 -526
rect 993 -538 997 -526
rect 1003 -538 1007 -526
rect 1021 -538 1025 -526
rect 936 -544 940 -538
rect 944 -544 948 -538
rect 64 -644 68 -634
rect 72 -644 76 -634
rect 100 -644 104 -634
rect 108 -644 112 -634
rect 116 -644 120 -634
rect 144 -644 148 -634
rect 152 -644 156 -634
rect 160 -644 164 -634
rect 195 -644 199 -634
rect 203 -644 207 -634
rect 264 -638 268 -628
rect 272 -638 276 -628
rect 300 -638 304 -628
rect 308 -638 312 -628
rect 316 -638 320 -628
rect 344 -638 348 -628
rect 352 -638 356 -628
rect 360 -638 364 -628
rect 395 -638 399 -628
rect 403 -638 407 -628
rect 450 -629 454 -616
rect 468 -629 472 -616
rect 492 -618 496 -611
rect 500 -618 504 -611
rect 885 -615 889 -609
rect 893 -615 897 -609
rect 450 -703 454 -690
rect 468 -703 472 -690
rect 492 -692 496 -685
rect 500 -692 504 -685
rect 63 -741 67 -731
rect 71 -741 75 -731
rect 99 -741 103 -731
rect 107 -741 111 -731
rect 115 -741 119 -731
rect 143 -741 147 -731
rect 151 -741 155 -731
rect 159 -741 163 -731
rect 194 -741 198 -731
rect 202 -741 206 -731
rect 263 -735 267 -725
rect 271 -735 275 -725
rect 299 -735 303 -725
rect 307 -735 311 -725
rect 315 -735 319 -725
rect 343 -735 347 -725
rect 351 -735 355 -725
rect 359 -735 363 -725
rect 394 -735 398 -725
rect 402 -735 406 -725
rect 450 -772 454 -759
rect 468 -772 472 -759
rect 492 -761 496 -754
rect 500 -761 504 -754
rect 64 -837 68 -827
rect 72 -837 76 -827
rect 100 -837 104 -827
rect 108 -837 112 -827
rect 116 -837 120 -827
rect 144 -837 148 -827
rect 152 -837 156 -827
rect 160 -837 164 -827
rect 195 -837 199 -827
rect 203 -837 207 -827
rect 264 -831 268 -821
rect 272 -831 276 -821
rect 300 -831 304 -821
rect 308 -831 312 -821
rect 316 -831 320 -821
rect 344 -831 348 -821
rect 352 -831 356 -821
rect 360 -831 364 -821
rect 395 -831 399 -821
rect 403 -831 407 -821
rect 450 -846 454 -833
rect 468 -846 472 -833
rect 492 -835 496 -828
rect 500 -835 504 -828
rect 548 -847 552 -623
rect 563 -847 568 -623
rect 602 -846 606 -622
rect 610 -846 614 -622
rect 635 -846 639 -622
rect 643 -846 647 -622
rect 666 -846 670 -622
rect 674 -846 678 -622
rect 700 -845 704 -621
rect 708 -845 712 -621
rect 721 -845 725 -621
rect 729 -845 733 -621
rect 738 -845 742 -621
rect 746 -845 750 -621
rect 756 -844 760 -620
rect 764 -844 768 -620
rect 801 -641 805 -634
rect 809 -641 813 -634
rect 924 -664 928 -652
rect 942 -664 946 -652
rect 952 -664 956 -652
rect 970 -664 974 -652
rect 1039 -660 1043 -650
rect 1047 -660 1051 -650
rect 1075 -660 1079 -650
rect 1083 -660 1087 -650
rect 1091 -660 1095 -650
rect 1119 -660 1123 -650
rect 1127 -660 1131 -650
rect 1135 -660 1139 -650
rect 1170 -660 1174 -650
rect 1178 -660 1182 -650
rect 885 -670 889 -664
rect 893 -670 897 -664
rect 802 -726 806 -719
rect 810 -726 814 -719
rect 896 -751 900 -745
rect 904 -751 908 -745
rect 935 -800 939 -788
rect 953 -800 957 -788
rect 963 -800 967 -788
rect 981 -800 985 -788
rect 896 -806 900 -800
rect 904 -806 908 -800
rect 1052 -802 1056 -792
rect 1060 -802 1064 -792
rect 1088 -802 1092 -792
rect 1096 -802 1100 -792
rect 1104 -802 1108 -792
rect 1132 -802 1136 -792
rect 1140 -802 1144 -792
rect 1148 -802 1152 -792
rect 1183 -802 1187 -792
rect 1191 -802 1195 -792
rect 805 -837 809 -830
rect 813 -837 817 -830
rect 905 -885 909 -879
rect 913 -885 917 -879
rect 806 -909 810 -902
rect 814 -909 818 -902
rect 266 -932 270 -922
rect 274 -932 278 -922
rect 302 -932 306 -922
rect 310 -932 314 -922
rect 318 -932 322 -922
rect 346 -932 350 -922
rect 354 -932 358 -922
rect 362 -932 366 -922
rect 397 -932 401 -922
rect 405 -932 409 -922
rect 944 -934 948 -922
rect 962 -934 966 -922
rect 972 -934 976 -922
rect 990 -934 994 -922
rect 1062 -925 1066 -915
rect 1070 -925 1074 -915
rect 1098 -925 1102 -915
rect 1106 -925 1110 -915
rect 1114 -925 1118 -915
rect 1142 -925 1146 -915
rect 1150 -925 1154 -915
rect 1158 -925 1162 -915
rect 1193 -925 1197 -915
rect 1201 -925 1205 -915
rect 905 -940 909 -934
rect 913 -940 917 -934
rect 631 -1001 635 -991
rect 639 -1001 643 -991
rect 667 -1001 671 -991
rect 675 -1001 679 -991
rect 683 -1001 687 -991
rect 711 -1001 715 -991
rect 719 -1001 723 -991
rect 727 -1001 731 -991
rect 762 -1001 766 -991
rect 770 -1001 774 -991
rect 910 -1034 914 -1028
rect 918 -1034 922 -1028
rect 949 -1083 953 -1071
rect 967 -1083 971 -1071
rect 977 -1083 981 -1071
rect 995 -1083 999 -1071
rect 1067 -1072 1071 -1062
rect 1075 -1072 1079 -1062
rect 1103 -1072 1107 -1062
rect 1111 -1072 1115 -1062
rect 1119 -1072 1123 -1062
rect 1147 -1072 1151 -1062
rect 1155 -1072 1159 -1062
rect 1163 -1072 1167 -1062
rect 1198 -1072 1202 -1062
rect 1206 -1072 1210 -1062
rect 910 -1089 914 -1083
rect 918 -1089 922 -1083
<< pdcontact >>
rect 523 -468 527 -456
rect 531 -468 535 -456
rect 71 -511 75 -486
rect 79 -511 83 -486
rect 87 -511 91 -486
rect 109 -511 113 -486
rect 117 -511 121 -486
rect 153 -511 157 -486
rect 161 -511 165 -486
rect 198 -511 202 -486
rect 206 -511 210 -486
rect 266 -508 270 -483
rect 274 -508 278 -483
rect 282 -508 286 -483
rect 304 -508 308 -483
rect 312 -508 316 -483
rect 348 -508 352 -483
rect 356 -508 360 -483
rect 393 -508 397 -483
rect 401 -508 405 -483
rect 562 -484 566 -460
rect 571 -484 575 -460
rect 580 -484 584 -460
rect 590 -490 594 -466
rect 599 -490 603 -466
rect 608 -490 612 -466
rect 663 -468 667 -456
rect 671 -468 675 -456
rect 702 -484 706 -460
rect 711 -484 715 -460
rect 720 -484 724 -460
rect 523 -523 527 -511
rect 531 -523 535 -511
rect 730 -490 734 -466
rect 739 -490 743 -466
rect 748 -490 752 -466
rect 798 -468 802 -456
rect 806 -468 810 -456
rect 837 -484 841 -460
rect 846 -484 850 -460
rect 855 -484 859 -460
rect 663 -523 667 -511
rect 671 -523 675 -511
rect 865 -490 869 -466
rect 874 -490 878 -466
rect 883 -490 887 -466
rect 936 -469 940 -457
rect 944 -469 948 -457
rect 975 -485 979 -461
rect 984 -485 988 -461
rect 993 -485 997 -461
rect 798 -523 802 -511
rect 806 -523 810 -511
rect 1003 -491 1007 -467
rect 1012 -491 1016 -467
rect 1021 -491 1025 -467
rect 936 -524 940 -512
rect 944 -524 948 -512
rect 68 -612 72 -587
rect 76 -612 80 -587
rect 84 -612 88 -587
rect 106 -612 110 -587
rect 114 -612 118 -587
rect 150 -612 154 -587
rect 158 -612 162 -587
rect 195 -612 199 -587
rect 203 -612 207 -587
rect 268 -606 272 -581
rect 276 -606 280 -581
rect 284 -606 288 -581
rect 306 -606 310 -581
rect 314 -606 318 -581
rect 350 -606 354 -581
rect 358 -606 362 -581
rect 395 -606 399 -581
rect 403 -606 407 -581
rect 450 -593 454 -581
rect 459 -593 463 -581
rect 468 -593 472 -581
rect 492 -593 496 -581
rect 500 -593 504 -581
rect 555 -591 559 -579
rect 563 -591 567 -579
rect 591 -591 595 -579
rect 599 -591 603 -579
rect 632 -591 636 -579
rect 640 -591 644 -579
rect 667 -591 671 -579
rect 675 -591 679 -579
rect 885 -595 889 -583
rect 893 -595 897 -583
rect 801 -616 805 -604
rect 809 -616 813 -604
rect 924 -611 928 -587
rect 933 -611 937 -587
rect 942 -611 946 -587
rect 450 -667 454 -655
rect 459 -667 463 -655
rect 468 -667 472 -655
rect 492 -667 496 -655
rect 500 -667 504 -655
rect 67 -709 71 -684
rect 75 -709 79 -684
rect 83 -709 87 -684
rect 105 -709 109 -684
rect 113 -709 117 -684
rect 149 -709 153 -684
rect 157 -709 161 -684
rect 194 -709 198 -684
rect 202 -709 206 -684
rect 267 -703 271 -678
rect 275 -703 279 -678
rect 283 -703 287 -678
rect 305 -703 309 -678
rect 313 -703 317 -678
rect 349 -703 353 -678
rect 357 -703 361 -678
rect 394 -703 398 -678
rect 402 -703 406 -678
rect 450 -736 454 -724
rect 459 -736 463 -724
rect 468 -736 472 -724
rect 492 -736 496 -724
rect 500 -736 504 -724
rect 68 -805 72 -780
rect 76 -805 80 -780
rect 84 -805 88 -780
rect 106 -805 110 -780
rect 114 -805 118 -780
rect 150 -805 154 -780
rect 158 -805 162 -780
rect 195 -805 199 -780
rect 203 -805 207 -780
rect 268 -799 272 -774
rect 276 -799 280 -774
rect 284 -799 288 -774
rect 306 -799 310 -774
rect 314 -799 318 -774
rect 350 -799 354 -774
rect 358 -799 362 -774
rect 395 -799 399 -774
rect 403 -799 407 -774
rect 450 -810 454 -798
rect 459 -810 463 -798
rect 468 -810 472 -798
rect 492 -810 496 -798
rect 500 -810 504 -798
rect 952 -617 956 -593
rect 961 -617 965 -593
rect 970 -617 974 -593
rect 885 -650 889 -638
rect 893 -650 897 -638
rect 1043 -628 1047 -603
rect 1051 -628 1055 -603
rect 1059 -628 1063 -603
rect 1081 -628 1085 -603
rect 1089 -628 1093 -603
rect 1125 -628 1129 -603
rect 1133 -628 1137 -603
rect 1170 -628 1174 -603
rect 1178 -628 1182 -603
rect 802 -701 806 -689
rect 810 -701 814 -689
rect 896 -731 900 -719
rect 904 -731 908 -719
rect 935 -747 939 -723
rect 944 -747 948 -723
rect 953 -747 957 -723
rect 963 -753 967 -729
rect 972 -753 976 -729
rect 981 -753 985 -729
rect 896 -786 900 -774
rect 904 -786 908 -774
rect 1056 -770 1060 -745
rect 1064 -770 1068 -745
rect 1072 -770 1076 -745
rect 1094 -770 1098 -745
rect 1102 -770 1106 -745
rect 1138 -770 1142 -745
rect 1146 -770 1150 -745
rect 1183 -770 1187 -745
rect 1191 -770 1195 -745
rect 805 -812 809 -800
rect 813 -812 817 -800
rect 905 -865 909 -853
rect 913 -865 917 -853
rect 270 -900 274 -875
rect 278 -900 282 -875
rect 286 -900 290 -875
rect 308 -900 312 -875
rect 316 -900 320 -875
rect 352 -900 356 -875
rect 360 -900 364 -875
rect 397 -900 401 -875
rect 405 -900 409 -875
rect 806 -884 810 -872
rect 814 -884 818 -872
rect 944 -881 948 -857
rect 953 -881 957 -857
rect 962 -881 966 -857
rect 972 -887 976 -863
rect 981 -887 985 -863
rect 990 -887 994 -863
rect 905 -920 909 -908
rect 913 -920 917 -908
rect 1066 -893 1070 -868
rect 1074 -893 1078 -868
rect 1082 -893 1086 -868
rect 1104 -893 1108 -868
rect 1112 -893 1116 -868
rect 1148 -893 1152 -868
rect 1156 -893 1160 -868
rect 1193 -893 1197 -868
rect 1201 -893 1205 -868
rect 635 -969 639 -944
rect 643 -969 647 -944
rect 651 -969 655 -944
rect 673 -969 677 -944
rect 681 -969 685 -944
rect 717 -969 721 -944
rect 725 -969 729 -944
rect 762 -969 766 -944
rect 770 -969 774 -944
rect 910 -1014 914 -1002
rect 918 -1014 922 -1002
rect 949 -1030 953 -1006
rect 958 -1030 962 -1006
rect 967 -1030 971 -1006
rect 977 -1036 981 -1012
rect 986 -1036 990 -1012
rect 995 -1036 999 -1012
rect 910 -1069 914 -1057
rect 918 -1069 922 -1057
rect 1071 -1040 1075 -1015
rect 1079 -1040 1083 -1015
rect 1087 -1040 1091 -1015
rect 1109 -1040 1113 -1015
rect 1117 -1040 1121 -1015
rect 1153 -1040 1157 -1015
rect 1161 -1040 1165 -1015
rect 1198 -1040 1202 -1015
rect 1206 -1040 1210 -1015
<< polysilicon >>
rect 528 -456 530 -453
rect 668 -456 670 -453
rect 803 -456 805 -453
rect 567 -460 569 -457
rect 577 -460 579 -457
rect 271 -483 273 -480
rect 279 -483 281 -480
rect 309 -483 311 -480
rect 353 -483 355 -480
rect 398 -483 400 -480
rect 528 -482 530 -468
rect 76 -486 78 -483
rect 84 -486 86 -483
rect 114 -486 116 -483
rect 158 -486 160 -483
rect 203 -486 205 -483
rect 595 -466 597 -463
rect 605 -466 607 -463
rect 528 -491 530 -488
rect 567 -493 569 -484
rect 577 -494 579 -484
rect 707 -460 709 -457
rect 717 -460 719 -457
rect 668 -482 670 -468
rect 735 -466 737 -463
rect 745 -466 747 -463
rect 76 -518 78 -511
rect 71 -522 78 -518
rect 72 -533 74 -522
rect 84 -530 86 -511
rect 114 -519 116 -511
rect 158 -519 160 -511
rect 108 -521 116 -519
rect 152 -521 160 -519
rect 108 -533 110 -521
rect 116 -533 118 -524
rect 152 -533 154 -521
rect 160 -533 162 -524
rect 203 -533 205 -511
rect 271 -515 273 -508
rect 266 -519 273 -515
rect 267 -530 269 -519
rect 279 -527 281 -508
rect 309 -516 311 -508
rect 353 -516 355 -508
rect 303 -518 311 -516
rect 347 -518 355 -516
rect 303 -530 305 -518
rect 311 -530 313 -521
rect 347 -530 349 -518
rect 355 -530 357 -521
rect 398 -530 400 -508
rect 528 -511 530 -508
rect 528 -537 530 -523
rect 567 -525 569 -498
rect 577 -525 579 -499
rect 595 -501 597 -490
rect 595 -525 597 -505
rect 605 -512 607 -490
rect 668 -491 670 -488
rect 707 -493 709 -484
rect 717 -494 719 -484
rect 941 -457 943 -454
rect 842 -460 844 -457
rect 852 -460 854 -457
rect 803 -482 805 -468
rect 870 -466 872 -463
rect 880 -466 882 -463
rect 668 -511 670 -508
rect 605 -525 607 -516
rect 668 -537 670 -523
rect 707 -525 709 -498
rect 717 -525 719 -499
rect 735 -501 737 -490
rect 735 -525 737 -505
rect 745 -512 747 -490
rect 803 -491 805 -488
rect 842 -493 844 -484
rect 852 -494 854 -484
rect 980 -461 982 -458
rect 990 -461 992 -458
rect 941 -483 943 -469
rect 1008 -467 1010 -464
rect 1018 -467 1020 -464
rect 803 -511 805 -508
rect 745 -525 747 -516
rect 803 -537 805 -523
rect 842 -525 844 -498
rect 852 -525 854 -499
rect 870 -501 872 -490
rect 870 -525 872 -505
rect 880 -512 882 -490
rect 941 -492 943 -489
rect 980 -494 982 -485
rect 990 -495 992 -485
rect 941 -512 943 -509
rect 880 -525 882 -516
rect 267 -543 269 -540
rect 303 -543 305 -540
rect 311 -543 313 -540
rect 347 -543 349 -540
rect 355 -543 357 -540
rect 398 -543 400 -540
rect 567 -540 569 -537
rect 577 -540 579 -537
rect 595 -540 597 -537
rect 605 -540 607 -537
rect 707 -540 709 -537
rect 717 -540 719 -537
rect 735 -540 737 -537
rect 745 -540 747 -537
rect 842 -540 844 -537
rect 852 -540 854 -537
rect 870 -540 872 -537
rect 880 -540 882 -537
rect 941 -538 943 -524
rect 980 -526 982 -499
rect 990 -526 992 -500
rect 1008 -502 1010 -491
rect 1008 -526 1010 -506
rect 1018 -513 1020 -491
rect 1018 -526 1020 -517
rect 72 -546 74 -543
rect 108 -546 110 -543
rect 116 -546 118 -543
rect 152 -546 154 -543
rect 160 -546 162 -543
rect 203 -546 205 -543
rect 528 -546 530 -543
rect 668 -546 670 -543
rect 803 -546 805 -543
rect 980 -541 982 -538
rect 990 -541 992 -538
rect 1008 -541 1010 -538
rect 1018 -541 1020 -538
rect 941 -547 943 -544
rect 273 -581 275 -578
rect 281 -581 283 -578
rect 311 -581 313 -578
rect 355 -581 357 -578
rect 400 -581 402 -578
rect 455 -581 457 -578
rect 465 -581 467 -578
rect 497 -581 499 -578
rect 560 -579 562 -576
rect 596 -579 598 -576
rect 637 -579 639 -576
rect 672 -579 674 -576
rect 73 -587 75 -584
rect 81 -587 83 -584
rect 111 -587 113 -584
rect 155 -587 157 -584
rect 200 -587 202 -584
rect 890 -583 892 -580
rect 73 -619 75 -612
rect 68 -623 75 -619
rect 69 -634 71 -623
rect 81 -631 83 -612
rect 111 -620 113 -612
rect 155 -620 157 -612
rect 105 -622 113 -620
rect 149 -622 157 -620
rect 105 -634 107 -622
rect 113 -634 115 -625
rect 149 -634 151 -622
rect 157 -634 159 -625
rect 200 -634 202 -612
rect 273 -613 275 -606
rect 268 -617 275 -613
rect 269 -628 271 -617
rect 281 -625 283 -606
rect 311 -614 313 -606
rect 355 -614 357 -606
rect 305 -616 313 -614
rect 349 -616 357 -614
rect 305 -628 307 -616
rect 313 -628 315 -619
rect 349 -628 351 -616
rect 357 -628 359 -619
rect 400 -628 402 -606
rect 455 -616 457 -593
rect 465 -616 467 -593
rect 497 -611 499 -593
rect 560 -606 562 -591
rect 596 -606 598 -591
rect 637 -606 639 -591
rect 672 -606 674 -591
rect 929 -587 931 -584
rect 939 -587 941 -584
rect 806 -604 808 -601
rect 497 -621 499 -618
rect 553 -623 555 -615
rect 560 -623 562 -615
rect 607 -622 609 -615
rect 640 -622 642 -615
rect 671 -622 673 -615
rect 705 -621 707 -614
rect 726 -621 728 -614
rect 743 -621 745 -614
rect 761 -620 763 -613
rect 890 -609 892 -595
rect 957 -593 959 -590
rect 967 -593 969 -590
rect 455 -633 457 -629
rect 465 -633 467 -629
rect 269 -641 271 -638
rect 305 -641 307 -638
rect 313 -641 315 -638
rect 349 -641 351 -638
rect 357 -641 359 -638
rect 400 -641 402 -638
rect 69 -647 71 -644
rect 105 -647 107 -644
rect 113 -647 115 -644
rect 149 -647 151 -644
rect 157 -647 159 -644
rect 200 -647 202 -644
rect 455 -655 457 -652
rect 465 -655 467 -652
rect 497 -655 499 -652
rect 272 -678 274 -675
rect 280 -678 282 -675
rect 310 -678 312 -675
rect 354 -678 356 -675
rect 399 -678 401 -675
rect 72 -684 74 -681
rect 80 -684 82 -681
rect 110 -684 112 -681
rect 154 -684 156 -681
rect 199 -684 201 -681
rect 455 -690 457 -667
rect 465 -690 467 -667
rect 497 -685 499 -667
rect 497 -695 499 -692
rect 72 -716 74 -709
rect 67 -720 74 -716
rect 68 -731 70 -720
rect 80 -728 82 -709
rect 110 -717 112 -709
rect 154 -717 156 -709
rect 104 -719 112 -717
rect 148 -719 156 -717
rect 104 -731 106 -719
rect 112 -731 114 -722
rect 148 -731 150 -719
rect 156 -731 158 -722
rect 199 -731 201 -709
rect 272 -710 274 -703
rect 267 -714 274 -710
rect 268 -725 270 -714
rect 280 -722 282 -703
rect 310 -711 312 -703
rect 354 -711 356 -703
rect 304 -713 312 -711
rect 348 -713 356 -711
rect 304 -725 306 -713
rect 312 -725 314 -716
rect 348 -725 350 -713
rect 356 -725 358 -716
rect 399 -725 401 -703
rect 455 -707 457 -703
rect 465 -707 467 -703
rect 455 -724 457 -721
rect 465 -724 467 -721
rect 497 -724 499 -721
rect 268 -738 270 -735
rect 304 -738 306 -735
rect 312 -738 314 -735
rect 348 -738 350 -735
rect 356 -738 358 -735
rect 399 -738 401 -735
rect 68 -744 70 -741
rect 104 -744 106 -741
rect 112 -744 114 -741
rect 148 -744 150 -741
rect 156 -744 158 -741
rect 199 -744 201 -741
rect 455 -759 457 -736
rect 465 -759 467 -736
rect 497 -754 499 -736
rect 273 -774 275 -771
rect 281 -774 283 -771
rect 311 -774 313 -771
rect 355 -774 357 -771
rect 400 -774 402 -771
rect 497 -764 499 -761
rect 73 -780 75 -777
rect 81 -780 83 -777
rect 111 -780 113 -777
rect 155 -780 157 -777
rect 200 -780 202 -777
rect 455 -776 457 -772
rect 465 -776 467 -772
rect 455 -798 457 -795
rect 465 -798 467 -795
rect 497 -798 499 -795
rect 73 -812 75 -805
rect 68 -816 75 -812
rect 69 -827 71 -816
rect 81 -824 83 -805
rect 111 -813 113 -805
rect 155 -813 157 -805
rect 105 -815 113 -813
rect 149 -815 157 -813
rect 105 -827 107 -815
rect 113 -827 115 -818
rect 149 -827 151 -815
rect 157 -827 159 -818
rect 200 -827 202 -805
rect 273 -806 275 -799
rect 268 -810 275 -806
rect 269 -821 271 -810
rect 281 -818 283 -799
rect 311 -807 313 -799
rect 355 -807 357 -799
rect 305 -809 313 -807
rect 349 -809 357 -807
rect 305 -821 307 -809
rect 313 -821 315 -812
rect 349 -821 351 -809
rect 357 -821 359 -812
rect 400 -821 402 -799
rect 269 -834 271 -831
rect 305 -834 307 -831
rect 313 -834 315 -831
rect 349 -834 351 -831
rect 357 -834 359 -831
rect 400 -834 402 -831
rect 455 -833 457 -810
rect 465 -833 467 -810
rect 497 -828 499 -810
rect 69 -840 71 -837
rect 105 -840 107 -837
rect 113 -840 115 -837
rect 149 -840 151 -837
rect 157 -840 159 -837
rect 200 -840 202 -837
rect 497 -838 499 -835
rect 455 -850 457 -846
rect 465 -850 467 -846
rect 806 -634 808 -616
rect 890 -618 892 -615
rect 929 -620 931 -611
rect 939 -621 941 -611
rect 1048 -603 1050 -600
rect 1056 -603 1058 -600
rect 1086 -603 1088 -600
rect 1130 -603 1132 -600
rect 1175 -603 1177 -600
rect 890 -638 892 -635
rect 806 -644 808 -641
rect 890 -664 892 -650
rect 929 -652 931 -625
rect 939 -652 941 -626
rect 957 -628 959 -617
rect 957 -652 959 -632
rect 967 -639 969 -617
rect 1048 -635 1050 -628
rect 1043 -639 1050 -635
rect 967 -652 969 -643
rect 1044 -650 1046 -639
rect 1056 -647 1058 -628
rect 1086 -636 1088 -628
rect 1130 -636 1132 -628
rect 1080 -638 1088 -636
rect 1124 -638 1132 -636
rect 1080 -650 1082 -638
rect 1088 -650 1090 -641
rect 1124 -650 1126 -638
rect 1132 -650 1134 -641
rect 1175 -650 1177 -628
rect 1044 -663 1046 -660
rect 1080 -663 1082 -660
rect 1088 -663 1090 -660
rect 1124 -663 1126 -660
rect 1132 -663 1134 -660
rect 1175 -663 1177 -660
rect 929 -667 931 -664
rect 939 -667 941 -664
rect 957 -667 959 -664
rect 967 -667 969 -664
rect 890 -673 892 -670
rect 807 -689 809 -686
rect 807 -719 809 -701
rect 901 -719 903 -716
rect 807 -729 809 -726
rect 940 -723 942 -720
rect 950 -723 952 -720
rect 901 -745 903 -731
rect 968 -729 970 -726
rect 978 -729 980 -726
rect 901 -754 903 -751
rect 940 -756 942 -747
rect 950 -757 952 -747
rect 1061 -745 1063 -742
rect 1069 -745 1071 -742
rect 1099 -745 1101 -742
rect 1143 -745 1145 -742
rect 1188 -745 1190 -742
rect 901 -774 903 -771
rect 810 -800 812 -797
rect 901 -800 903 -786
rect 940 -788 942 -761
rect 950 -788 952 -762
rect 968 -764 970 -753
rect 968 -788 970 -768
rect 978 -775 980 -753
rect 1061 -777 1063 -770
rect 978 -788 980 -779
rect 1056 -781 1063 -777
rect 1057 -792 1059 -781
rect 1069 -789 1071 -770
rect 1099 -778 1101 -770
rect 1143 -778 1145 -770
rect 1093 -780 1101 -778
rect 1137 -780 1145 -778
rect 1093 -792 1095 -780
rect 1101 -792 1103 -783
rect 1137 -792 1139 -780
rect 1145 -792 1147 -783
rect 1188 -792 1190 -770
rect 940 -803 942 -800
rect 950 -803 952 -800
rect 968 -803 970 -800
rect 978 -803 980 -800
rect 1057 -805 1059 -802
rect 1093 -805 1095 -802
rect 1101 -805 1103 -802
rect 1137 -805 1139 -802
rect 1145 -805 1147 -802
rect 1188 -805 1190 -802
rect 901 -809 903 -806
rect 810 -830 812 -812
rect 810 -840 812 -837
rect 553 -850 555 -847
rect 560 -850 562 -847
rect 607 -850 609 -846
rect 640 -850 642 -846
rect 671 -850 673 -846
rect 705 -849 707 -845
rect 726 -849 728 -845
rect 743 -849 745 -845
rect 761 -848 763 -844
rect 910 -853 912 -850
rect 949 -857 951 -854
rect 959 -857 961 -854
rect 811 -872 813 -869
rect 275 -875 277 -872
rect 283 -875 285 -872
rect 313 -875 315 -872
rect 357 -875 359 -872
rect 402 -875 404 -872
rect 910 -879 912 -865
rect 275 -907 277 -900
rect 270 -911 277 -907
rect 271 -922 273 -911
rect 283 -919 285 -900
rect 313 -908 315 -900
rect 357 -908 359 -900
rect 307 -910 315 -908
rect 351 -910 359 -908
rect 307 -922 309 -910
rect 315 -922 317 -913
rect 351 -922 353 -910
rect 359 -922 361 -913
rect 402 -922 404 -900
rect 811 -902 813 -884
rect 977 -863 979 -860
rect 987 -863 989 -860
rect 910 -888 912 -885
rect 949 -890 951 -881
rect 959 -891 961 -881
rect 1071 -868 1073 -865
rect 1079 -868 1081 -865
rect 1109 -868 1111 -865
rect 1153 -868 1155 -865
rect 1198 -868 1200 -865
rect 910 -908 912 -905
rect 811 -912 813 -909
rect 271 -935 273 -932
rect 307 -935 309 -932
rect 315 -935 317 -932
rect 351 -935 353 -932
rect 359 -935 361 -932
rect 402 -935 404 -932
rect 910 -934 912 -920
rect 949 -922 951 -895
rect 959 -922 961 -896
rect 977 -898 979 -887
rect 977 -922 979 -902
rect 987 -909 989 -887
rect 1071 -900 1073 -893
rect 1066 -904 1073 -900
rect 987 -922 989 -913
rect 1067 -915 1069 -904
rect 1079 -912 1081 -893
rect 1109 -901 1111 -893
rect 1153 -901 1155 -893
rect 1103 -903 1111 -901
rect 1147 -903 1155 -901
rect 1103 -915 1105 -903
rect 1111 -915 1113 -906
rect 1147 -915 1149 -903
rect 1155 -915 1157 -906
rect 1198 -915 1200 -893
rect 1067 -928 1069 -925
rect 1103 -928 1105 -925
rect 1111 -928 1113 -925
rect 1147 -928 1149 -925
rect 1155 -928 1157 -925
rect 1198 -928 1200 -925
rect 949 -937 951 -934
rect 959 -937 961 -934
rect 977 -937 979 -934
rect 987 -937 989 -934
rect 640 -944 642 -941
rect 648 -944 650 -941
rect 678 -944 680 -941
rect 722 -944 724 -941
rect 767 -944 769 -941
rect 910 -943 912 -940
rect 640 -976 642 -969
rect 635 -980 642 -976
rect 636 -991 638 -980
rect 648 -988 650 -969
rect 678 -977 680 -969
rect 722 -977 724 -969
rect 672 -979 680 -977
rect 716 -979 724 -977
rect 672 -991 674 -979
rect 680 -991 682 -982
rect 716 -991 718 -979
rect 724 -991 726 -982
rect 767 -991 769 -969
rect 636 -1004 638 -1001
rect 672 -1004 674 -1001
rect 680 -1004 682 -1001
rect 716 -1004 718 -1001
rect 724 -1004 726 -1001
rect 767 -1004 769 -1001
rect 915 -1002 917 -999
rect 954 -1006 956 -1003
rect 964 -1006 966 -1003
rect 915 -1028 917 -1014
rect 982 -1012 984 -1009
rect 992 -1012 994 -1009
rect 915 -1037 917 -1034
rect 954 -1039 956 -1030
rect 964 -1040 966 -1030
rect 1076 -1015 1078 -1012
rect 1084 -1015 1086 -1012
rect 1114 -1015 1116 -1012
rect 1158 -1015 1160 -1012
rect 1203 -1015 1205 -1012
rect 915 -1057 917 -1054
rect 915 -1083 917 -1069
rect 954 -1071 956 -1044
rect 964 -1071 966 -1045
rect 982 -1047 984 -1036
rect 982 -1071 984 -1051
rect 992 -1058 994 -1036
rect 1076 -1047 1078 -1040
rect 1071 -1051 1078 -1047
rect 1072 -1062 1074 -1051
rect 1084 -1059 1086 -1040
rect 1114 -1048 1116 -1040
rect 1158 -1048 1160 -1040
rect 1108 -1050 1116 -1048
rect 1152 -1050 1160 -1048
rect 1108 -1062 1110 -1050
rect 1116 -1062 1118 -1053
rect 1152 -1062 1154 -1050
rect 1160 -1062 1162 -1053
rect 1203 -1062 1205 -1040
rect 992 -1071 994 -1062
rect 1072 -1075 1074 -1072
rect 1108 -1075 1110 -1072
rect 1116 -1075 1118 -1072
rect 1152 -1075 1154 -1072
rect 1160 -1075 1162 -1072
rect 1203 -1075 1205 -1072
rect 954 -1086 956 -1083
rect 964 -1086 966 -1083
rect 982 -1086 984 -1083
rect 992 -1086 994 -1083
rect 915 -1092 917 -1089
<< polycontact >>
rect 524 -479 528 -475
rect 664 -479 668 -475
rect 67 -522 71 -518
rect 80 -530 84 -526
rect 91 -522 95 -518
rect 103 -530 108 -525
rect 118 -530 122 -526
rect 147 -530 152 -525
rect 199 -525 203 -520
rect 162 -530 166 -526
rect 262 -519 266 -515
rect 275 -527 279 -523
rect 286 -519 290 -515
rect 298 -527 303 -522
rect 313 -527 317 -523
rect 342 -527 347 -522
rect 394 -522 398 -517
rect 357 -527 361 -523
rect 524 -534 528 -530
rect 593 -505 597 -501
rect 799 -479 803 -475
rect 604 -516 608 -512
rect 664 -534 668 -530
rect 733 -505 737 -501
rect 937 -480 941 -476
rect 744 -516 748 -512
rect 799 -534 803 -530
rect 868 -505 872 -501
rect 879 -516 883 -512
rect 937 -535 941 -531
rect 1006 -506 1010 -502
rect 1017 -517 1021 -513
rect 451 -606 455 -602
rect 64 -623 68 -619
rect 77 -631 81 -627
rect 88 -623 92 -619
rect 100 -631 105 -626
rect 115 -631 119 -627
rect 144 -631 149 -626
rect 196 -626 200 -621
rect 159 -631 163 -627
rect 264 -617 268 -613
rect 277 -625 281 -621
rect 288 -617 292 -613
rect 300 -625 305 -620
rect 315 -625 319 -621
rect 344 -625 349 -620
rect 396 -620 400 -615
rect 359 -625 363 -621
rect 461 -613 465 -609
rect 493 -607 497 -603
rect 556 -606 560 -602
rect 592 -606 596 -602
rect 633 -606 637 -602
rect 668 -606 672 -602
rect 549 -619 553 -615
rect 562 -619 566 -615
rect 603 -619 607 -615
rect 636 -619 640 -615
rect 667 -619 671 -615
rect 701 -618 705 -614
rect 722 -618 726 -614
rect 739 -618 743 -614
rect 757 -617 761 -613
rect 886 -606 890 -602
rect 451 -680 455 -676
rect 461 -687 465 -683
rect 493 -681 497 -677
rect 63 -720 67 -716
rect 76 -728 80 -724
rect 87 -720 91 -716
rect 99 -728 104 -723
rect 114 -728 118 -724
rect 143 -728 148 -723
rect 195 -723 199 -718
rect 158 -728 162 -724
rect 263 -714 267 -710
rect 276 -722 280 -718
rect 287 -714 291 -710
rect 299 -722 304 -717
rect 314 -722 318 -718
rect 343 -722 348 -717
rect 395 -717 399 -712
rect 358 -722 362 -718
rect 451 -749 455 -745
rect 461 -756 465 -752
rect 493 -750 497 -746
rect 64 -816 68 -812
rect 77 -824 81 -820
rect 88 -816 92 -812
rect 100 -824 105 -819
rect 115 -824 119 -820
rect 144 -824 149 -819
rect 196 -819 200 -814
rect 159 -824 163 -820
rect 264 -810 268 -806
rect 277 -818 281 -814
rect 288 -810 292 -806
rect 300 -818 305 -813
rect 315 -818 319 -814
rect 344 -818 349 -813
rect 396 -813 400 -808
rect 359 -818 363 -814
rect 451 -823 455 -819
rect 461 -830 465 -826
rect 493 -824 497 -820
rect 802 -630 806 -626
rect 886 -661 890 -657
rect 955 -632 959 -628
rect 1039 -639 1043 -635
rect 966 -643 970 -639
rect 1052 -647 1056 -643
rect 1063 -639 1067 -635
rect 1075 -647 1080 -642
rect 1090 -647 1094 -643
rect 1119 -647 1124 -642
rect 1171 -642 1175 -637
rect 1134 -647 1138 -643
rect 803 -715 807 -711
rect 897 -742 901 -738
rect 897 -797 901 -793
rect 966 -768 970 -764
rect 977 -779 981 -775
rect 1052 -781 1056 -777
rect 1065 -789 1069 -785
rect 1076 -781 1080 -777
rect 1088 -789 1093 -784
rect 1103 -789 1107 -785
rect 1132 -789 1137 -784
rect 1184 -784 1188 -779
rect 1147 -789 1151 -785
rect 806 -826 810 -822
rect 906 -876 910 -872
rect 807 -898 811 -894
rect 266 -911 270 -907
rect 279 -919 283 -915
rect 290 -911 294 -907
rect 302 -919 307 -914
rect 317 -919 321 -915
rect 346 -919 351 -914
rect 398 -914 402 -909
rect 361 -919 365 -915
rect 906 -931 910 -927
rect 975 -902 979 -898
rect 1062 -904 1066 -900
rect 986 -913 990 -909
rect 1075 -912 1079 -908
rect 1086 -904 1090 -900
rect 1098 -912 1103 -907
rect 1113 -912 1117 -908
rect 1142 -912 1147 -907
rect 1194 -907 1198 -902
rect 1157 -912 1161 -908
rect 631 -980 635 -976
rect 644 -988 648 -984
rect 655 -980 659 -976
rect 667 -988 672 -983
rect 682 -988 686 -984
rect 711 -988 716 -983
rect 763 -983 767 -978
rect 726 -988 730 -984
rect 911 -1025 915 -1021
rect 911 -1080 915 -1076
rect 980 -1051 984 -1047
rect 1067 -1051 1071 -1047
rect 991 -1062 995 -1058
rect 1080 -1059 1084 -1055
rect 1091 -1051 1095 -1047
rect 1103 -1059 1108 -1054
rect 1118 -1059 1122 -1055
rect 1147 -1059 1152 -1054
rect 1199 -1054 1203 -1049
rect 1162 -1059 1166 -1055
<< metal1 >>
rect 522 -450 550 -447
rect 662 -450 690 -447
rect 797 -450 825 -447
rect 523 -456 526 -450
rect 547 -451 550 -450
rect 547 -454 618 -451
rect 65 -480 218 -476
rect 260 -477 413 -473
rect 71 -486 75 -480
rect 109 -486 113 -480
rect 153 -486 157 -480
rect 198 -486 202 -480
rect 266 -483 270 -477
rect 304 -483 308 -477
rect 348 -483 352 -477
rect 393 -483 397 -477
rect 506 -480 509 -477
rect 514 -479 524 -476
rect 532 -476 535 -468
rect 562 -460 565 -454
rect 581 -460 584 -454
rect 663 -456 666 -450
rect 687 -451 690 -450
rect 687 -454 758 -451
rect 532 -479 553 -476
rect 532 -482 535 -479
rect 121 -511 134 -486
rect 165 -511 178 -486
rect 316 -508 329 -483
rect 360 -508 373 -483
rect 523 -492 526 -488
rect 517 -494 541 -492
rect 517 -495 535 -494
rect 540 -495 541 -494
rect 550 -502 553 -479
rect 591 -460 611 -457
rect 591 -466 594 -460
rect 608 -466 611 -460
rect 572 -487 575 -484
rect 572 -490 590 -487
rect 646 -480 649 -477
rect 654 -479 664 -476
rect 672 -476 675 -468
rect 702 -460 705 -454
rect 721 -460 724 -454
rect 798 -456 801 -450
rect 822 -451 825 -450
rect 935 -451 963 -448
rect 822 -454 893 -451
rect 672 -479 693 -476
rect 672 -482 675 -479
rect 600 -497 603 -490
rect 663 -492 666 -488
rect 657 -494 681 -492
rect 657 -495 675 -494
rect 600 -500 617 -497
rect 522 -503 541 -502
rect 517 -505 541 -503
rect 550 -505 593 -502
rect 60 -522 67 -518
rect 71 -530 80 -526
rect 87 -533 91 -511
rect 95 -522 96 -518
rect 131 -520 134 -511
rect 175 -520 178 -511
rect 131 -525 143 -520
rect 175 -525 199 -520
rect 206 -521 210 -511
rect 255 -519 262 -515
rect 95 -527 103 -525
rect 100 -530 103 -527
rect 122 -530 123 -526
rect 131 -533 134 -525
rect 139 -530 147 -525
rect 166 -530 167 -526
rect 175 -533 178 -525
rect 206 -526 219 -521
rect 206 -533 210 -526
rect 266 -527 275 -523
rect 282 -530 286 -508
rect 290 -519 291 -515
rect 326 -517 329 -508
rect 370 -517 373 -508
rect 326 -522 338 -517
rect 370 -522 394 -517
rect 401 -518 405 -508
rect 523 -511 526 -505
rect 614 -511 617 -500
rect 680 -495 681 -494
rect 690 -502 693 -479
rect 731 -460 751 -457
rect 731 -466 734 -460
rect 748 -466 751 -460
rect 712 -487 715 -484
rect 712 -490 730 -487
rect 781 -480 784 -477
rect 789 -479 799 -476
rect 807 -476 810 -468
rect 837 -460 840 -454
rect 856 -460 859 -454
rect 936 -457 939 -451
rect 960 -452 963 -451
rect 960 -455 1031 -452
rect 807 -479 828 -476
rect 807 -482 810 -479
rect 740 -497 743 -490
rect 798 -492 801 -488
rect 792 -494 816 -492
rect 792 -495 810 -494
rect 740 -500 757 -497
rect 662 -503 681 -502
rect 657 -505 681 -503
rect 690 -505 733 -502
rect 663 -511 666 -505
rect 754 -511 757 -500
rect 815 -495 816 -494
rect 825 -502 828 -479
rect 866 -460 886 -457
rect 866 -466 869 -460
rect 883 -466 886 -460
rect 847 -487 850 -484
rect 847 -490 865 -487
rect 919 -481 922 -478
rect 927 -480 937 -477
rect 945 -477 948 -469
rect 975 -461 978 -455
rect 994 -461 997 -455
rect 945 -480 966 -477
rect 945 -483 948 -480
rect 875 -497 878 -490
rect 936 -493 939 -489
rect 930 -495 954 -493
rect 930 -496 948 -495
rect 875 -500 892 -497
rect 797 -503 816 -502
rect 792 -505 816 -503
rect 825 -505 868 -502
rect 798 -511 801 -505
rect 889 -511 892 -500
rect 953 -496 954 -495
rect 963 -503 966 -480
rect 1004 -461 1024 -458
rect 1004 -467 1007 -461
rect 1021 -467 1024 -461
rect 985 -488 988 -485
rect 985 -491 1003 -488
rect 1013 -498 1016 -491
rect 1013 -501 1030 -498
rect 935 -504 954 -503
rect 930 -506 954 -504
rect 963 -506 1006 -503
rect 290 -524 298 -522
rect 295 -527 298 -524
rect 317 -527 318 -523
rect 326 -530 329 -522
rect 334 -527 342 -522
rect 361 -527 362 -523
rect 370 -530 373 -522
rect 401 -523 414 -518
rect 579 -516 604 -513
rect 614 -515 627 -511
rect 579 -518 582 -516
rect 401 -530 405 -523
rect 79 -543 91 -533
rect 123 -543 134 -533
rect 167 -543 178 -533
rect 274 -540 286 -530
rect 318 -540 329 -530
rect 362 -540 373 -530
rect 506 -534 509 -531
rect 514 -534 524 -531
rect 532 -531 535 -523
rect 544 -521 582 -518
rect 614 -519 617 -515
rect 544 -531 547 -521
rect 585 -522 617 -519
rect 585 -525 588 -522
rect 532 -534 547 -531
rect 532 -537 535 -534
rect 67 -548 71 -543
rect 103 -548 107 -543
rect 147 -548 151 -543
rect 198 -548 202 -543
rect 262 -545 266 -540
rect 298 -545 302 -540
rect 342 -545 346 -540
rect 393 -545 397 -540
rect 584 -528 590 -525
rect 66 -552 210 -548
rect 261 -549 405 -545
rect 523 -547 526 -543
rect 544 -544 549 -541
rect 562 -541 565 -537
rect 609 -541 612 -537
rect 554 -544 618 -541
rect 544 -547 547 -544
rect 517 -550 547 -547
rect 623 -555 627 -515
rect 719 -516 744 -513
rect 754 -515 766 -511
rect 719 -518 722 -516
rect 646 -534 649 -531
rect 654 -534 664 -531
rect 672 -531 675 -523
rect 684 -521 722 -518
rect 754 -519 757 -515
rect 684 -531 687 -521
rect 725 -522 757 -519
rect 725 -525 728 -522
rect 672 -534 687 -531
rect 672 -537 675 -534
rect 724 -528 730 -525
rect 663 -547 666 -543
rect 684 -544 689 -541
rect 702 -541 705 -537
rect 749 -541 752 -537
rect 694 -544 758 -541
rect 684 -547 687 -544
rect 657 -550 687 -547
rect 762 -556 766 -515
rect 854 -516 879 -513
rect 889 -515 900 -511
rect 854 -518 857 -516
rect 781 -534 784 -531
rect 789 -534 799 -531
rect 807 -531 810 -523
rect 819 -521 857 -518
rect 889 -519 892 -515
rect 819 -531 822 -521
rect 860 -522 892 -519
rect 860 -525 863 -522
rect 807 -534 822 -531
rect 807 -537 810 -534
rect 859 -528 865 -525
rect 798 -547 801 -543
rect 819 -544 824 -541
rect 837 -541 840 -537
rect 884 -541 887 -537
rect 829 -544 893 -541
rect 819 -547 822 -544
rect 792 -550 822 -547
rect 896 -555 900 -515
rect 936 -512 939 -506
rect 1027 -512 1030 -501
rect 992 -517 1017 -514
rect 1027 -516 1042 -512
rect 992 -519 995 -517
rect 919 -535 922 -532
rect 927 -535 937 -532
rect 945 -532 948 -524
rect 957 -522 995 -519
rect 1027 -520 1030 -516
rect 957 -532 960 -522
rect 998 -523 1030 -520
rect 998 -526 1001 -523
rect 945 -535 960 -532
rect 945 -538 948 -535
rect 997 -529 1003 -526
rect 936 -548 939 -544
rect 957 -545 962 -542
rect 975 -542 978 -538
rect 1022 -542 1025 -538
rect 967 -545 1031 -542
rect 957 -548 960 -545
rect 930 -551 960 -548
rect 1038 -554 1042 -516
rect 762 -560 769 -556
rect 893 -559 900 -555
rect 262 -575 415 -571
rect 442 -575 513 -572
rect 548 -573 576 -570
rect 584 -573 612 -570
rect 625 -573 653 -570
rect 660 -573 688 -570
rect 62 -581 215 -577
rect 268 -581 272 -575
rect 306 -581 310 -575
rect 350 -581 354 -575
rect 395 -581 399 -575
rect 450 -581 454 -575
rect 468 -581 472 -575
rect 68 -587 72 -581
rect 106 -587 110 -581
rect 150 -587 154 -581
rect 195 -587 199 -581
rect 118 -612 131 -587
rect 162 -612 175 -587
rect 318 -606 331 -581
rect 362 -606 375 -581
rect 492 -581 495 -575
rect 555 -579 558 -573
rect 591 -579 594 -573
rect 632 -579 635 -573
rect 667 -579 670 -573
rect 884 -577 912 -574
rect 459 -596 462 -593
rect 459 -599 472 -596
rect 442 -606 451 -602
rect 469 -603 472 -599
rect 501 -603 504 -593
rect 57 -623 64 -619
rect 68 -631 77 -627
rect 84 -634 88 -612
rect 92 -623 93 -619
rect 128 -621 131 -612
rect 172 -621 175 -612
rect 128 -626 140 -621
rect 172 -626 196 -621
rect 203 -622 207 -612
rect 257 -617 264 -613
rect 92 -628 100 -626
rect 97 -631 100 -628
rect 119 -631 120 -627
rect 128 -634 131 -626
rect 136 -631 144 -626
rect 163 -631 164 -627
rect 172 -634 175 -626
rect 203 -627 216 -622
rect 268 -625 277 -621
rect 203 -634 207 -627
rect 284 -628 288 -606
rect 292 -617 293 -613
rect 328 -615 331 -606
rect 372 -615 375 -606
rect 328 -620 340 -615
rect 372 -620 396 -615
rect 403 -616 407 -606
rect 469 -607 493 -603
rect 501 -606 513 -603
rect 548 -606 556 -602
rect 564 -606 567 -591
rect 584 -606 592 -602
rect 600 -606 603 -591
rect 625 -606 633 -602
rect 641 -606 644 -591
rect 660 -606 668 -602
rect 676 -606 679 -591
rect 885 -583 888 -577
rect 909 -578 912 -577
rect 909 -581 980 -578
rect 790 -598 822 -595
rect 801 -604 804 -598
rect 442 -613 461 -609
rect 469 -616 472 -607
rect 501 -611 504 -606
rect 292 -622 300 -620
rect 297 -625 300 -622
rect 319 -625 320 -621
rect 328 -628 331 -620
rect 336 -625 344 -620
rect 363 -625 364 -621
rect 372 -628 375 -620
rect 403 -621 416 -616
rect 403 -628 407 -621
rect 76 -644 88 -634
rect 120 -644 131 -634
rect 164 -644 175 -634
rect 276 -638 288 -628
rect 320 -638 331 -628
rect 364 -638 375 -628
rect 450 -635 453 -629
rect 492 -635 495 -618
rect 546 -619 549 -615
rect 566 -619 572 -615
rect 600 -619 603 -615
rect 633 -619 636 -615
rect 664 -619 667 -615
rect 674 -622 678 -615
rect 698 -618 701 -614
rect 708 -621 712 -614
rect 719 -618 722 -614
rect 729 -621 733 -614
rect 736 -618 739 -614
rect 746 -621 750 -614
rect 754 -617 757 -613
rect 764 -620 768 -613
rect 868 -607 871 -604
rect 876 -606 886 -603
rect 894 -603 897 -595
rect 924 -587 927 -581
rect 943 -587 946 -581
rect 894 -606 915 -603
rect 894 -609 897 -606
rect 442 -638 495 -635
rect 264 -643 268 -638
rect 300 -643 304 -638
rect 344 -643 348 -638
rect 395 -643 399 -638
rect 64 -649 68 -644
rect 100 -649 104 -644
rect 144 -649 148 -644
rect 195 -649 199 -644
rect 263 -647 407 -643
rect 442 -649 513 -646
rect 63 -653 207 -649
rect 450 -655 454 -649
rect 468 -655 472 -649
rect 492 -655 495 -649
rect 261 -672 414 -668
rect 459 -670 462 -667
rect 61 -678 214 -674
rect 267 -678 271 -672
rect 305 -678 309 -672
rect 349 -678 353 -672
rect 394 -678 398 -672
rect 459 -673 472 -670
rect 67 -684 71 -678
rect 105 -684 109 -678
rect 149 -684 153 -678
rect 194 -684 198 -678
rect 117 -709 130 -684
rect 161 -709 174 -684
rect 317 -703 330 -678
rect 361 -703 374 -678
rect 442 -680 451 -676
rect 469 -677 472 -673
rect 501 -677 504 -667
rect 469 -681 493 -677
rect 501 -680 513 -677
rect 442 -687 461 -683
rect 469 -690 472 -681
rect 501 -685 504 -680
rect 56 -720 63 -716
rect 67 -728 76 -724
rect 83 -731 87 -709
rect 91 -720 92 -716
rect 127 -718 130 -709
rect 171 -718 174 -709
rect 127 -723 139 -718
rect 171 -723 195 -718
rect 202 -719 206 -709
rect 256 -714 263 -710
rect 91 -725 99 -723
rect 96 -728 99 -725
rect 118 -728 119 -724
rect 127 -731 130 -723
rect 135 -728 143 -723
rect 162 -728 163 -724
rect 171 -731 174 -723
rect 202 -724 215 -719
rect 267 -722 276 -718
rect 202 -731 206 -724
rect 283 -725 287 -703
rect 291 -714 292 -710
rect 327 -712 330 -703
rect 371 -712 374 -703
rect 327 -717 339 -712
rect 371 -717 395 -712
rect 402 -713 406 -703
rect 450 -709 453 -703
rect 492 -709 495 -692
rect 442 -712 495 -709
rect 291 -719 299 -717
rect 296 -722 299 -719
rect 318 -722 319 -718
rect 327 -725 330 -717
rect 335 -722 343 -717
rect 362 -722 363 -718
rect 371 -725 374 -717
rect 402 -718 415 -713
rect 442 -718 513 -715
rect 402 -725 406 -718
rect 75 -741 87 -731
rect 119 -741 130 -731
rect 163 -741 174 -731
rect 275 -735 287 -725
rect 319 -735 330 -725
rect 363 -735 374 -725
rect 450 -724 454 -718
rect 468 -724 472 -718
rect 263 -740 267 -735
rect 299 -740 303 -735
rect 343 -740 347 -735
rect 394 -740 398 -735
rect 492 -724 495 -718
rect 459 -739 462 -736
rect 63 -746 67 -741
rect 99 -746 103 -741
rect 143 -746 147 -741
rect 194 -746 198 -741
rect 262 -744 406 -740
rect 459 -742 472 -739
rect 62 -750 206 -746
rect 442 -749 451 -745
rect 469 -746 472 -742
rect 501 -746 504 -736
rect 469 -750 493 -746
rect 501 -749 513 -746
rect 442 -756 461 -752
rect 469 -759 472 -750
rect 501 -754 504 -749
rect 262 -768 415 -764
rect 62 -774 215 -770
rect 268 -774 272 -768
rect 306 -774 310 -768
rect 350 -774 354 -768
rect 395 -774 399 -768
rect 68 -780 72 -774
rect 106 -780 110 -774
rect 150 -780 154 -774
rect 195 -780 199 -774
rect 118 -805 131 -780
rect 162 -805 175 -780
rect 318 -799 331 -774
rect 362 -799 375 -774
rect 450 -778 453 -772
rect 492 -778 495 -761
rect 442 -781 495 -778
rect 442 -792 513 -789
rect 57 -816 64 -812
rect 68 -824 77 -820
rect 84 -827 88 -805
rect 92 -816 93 -812
rect 128 -814 131 -805
rect 172 -814 175 -805
rect 128 -819 140 -814
rect 172 -819 196 -814
rect 203 -815 207 -805
rect 257 -810 264 -806
rect 92 -821 100 -819
rect 97 -824 100 -821
rect 119 -824 120 -820
rect 128 -827 131 -819
rect 136 -824 144 -819
rect 163 -824 164 -820
rect 172 -827 175 -819
rect 203 -820 216 -815
rect 268 -818 277 -814
rect 203 -827 207 -820
rect 284 -821 288 -799
rect 292 -810 293 -806
rect 328 -808 331 -799
rect 372 -808 375 -799
rect 328 -813 340 -808
rect 372 -813 396 -808
rect 403 -809 407 -799
rect 450 -798 454 -792
rect 468 -798 472 -792
rect 292 -815 300 -813
rect 297 -818 300 -815
rect 319 -818 320 -814
rect 328 -821 331 -813
rect 336 -818 344 -813
rect 363 -818 364 -814
rect 372 -821 375 -813
rect 403 -814 416 -809
rect 492 -798 495 -792
rect 459 -813 462 -810
rect 403 -821 407 -814
rect 459 -816 472 -813
rect 76 -837 88 -827
rect 120 -837 131 -827
rect 164 -837 175 -827
rect 276 -831 288 -821
rect 320 -831 331 -821
rect 364 -831 375 -821
rect 442 -823 451 -819
rect 469 -820 472 -816
rect 501 -820 504 -810
rect 469 -824 493 -820
rect 501 -823 513 -820
rect 442 -830 461 -826
rect 264 -836 268 -831
rect 300 -836 304 -831
rect 344 -836 348 -831
rect 395 -836 399 -831
rect 469 -833 472 -824
rect 501 -828 504 -823
rect 64 -842 68 -837
rect 100 -842 104 -837
rect 144 -842 148 -837
rect 195 -842 199 -837
rect 263 -840 407 -836
rect 63 -846 207 -842
rect 450 -852 453 -846
rect 492 -852 495 -835
rect 442 -855 495 -852
rect 548 -856 552 -847
rect 563 -848 568 -847
rect 602 -848 606 -846
rect 563 -853 606 -848
rect 610 -848 614 -846
rect 635 -848 639 -846
rect 610 -853 639 -848
rect 643 -848 647 -846
rect 810 -626 813 -616
rect 885 -619 888 -615
rect 879 -621 903 -619
rect 879 -622 897 -621
rect 790 -630 802 -626
rect 810 -629 822 -626
rect 810 -634 813 -629
rect 902 -622 903 -621
rect 912 -629 915 -606
rect 953 -587 973 -584
rect 953 -593 956 -587
rect 970 -593 973 -587
rect 934 -614 937 -611
rect 934 -617 952 -614
rect 1037 -597 1190 -593
rect 1043 -603 1047 -597
rect 1081 -603 1085 -597
rect 1125 -603 1129 -597
rect 1170 -603 1174 -597
rect 962 -624 965 -617
rect 962 -627 979 -624
rect 884 -630 903 -629
rect 879 -632 903 -630
rect 912 -632 955 -629
rect 885 -638 888 -632
rect 976 -638 979 -627
rect 1093 -628 1106 -603
rect 1137 -628 1150 -603
rect 801 -658 804 -641
rect 941 -643 966 -640
rect 976 -642 989 -638
rect 1032 -639 1039 -635
rect 941 -645 944 -643
rect 790 -661 804 -658
rect 868 -661 871 -658
rect 876 -661 886 -658
rect 894 -658 897 -650
rect 906 -648 944 -645
rect 976 -646 979 -642
rect 906 -658 909 -648
rect 947 -649 979 -646
rect 947 -652 950 -649
rect 894 -661 909 -658
rect 894 -664 897 -661
rect 946 -655 952 -652
rect 885 -674 888 -670
rect 906 -671 911 -668
rect 924 -668 927 -664
rect 971 -668 974 -664
rect 916 -671 980 -668
rect 906 -674 909 -671
rect 879 -677 909 -674
rect 791 -683 823 -680
rect 985 -682 989 -642
rect 1043 -647 1052 -643
rect 1059 -650 1063 -628
rect 1067 -639 1068 -635
rect 1103 -637 1106 -628
rect 1147 -637 1150 -628
rect 1103 -642 1115 -637
rect 1147 -642 1171 -637
rect 1178 -638 1182 -628
rect 1067 -644 1075 -642
rect 1072 -647 1075 -644
rect 1094 -647 1095 -643
rect 1103 -650 1106 -642
rect 1111 -647 1119 -642
rect 1138 -647 1139 -643
rect 1147 -650 1150 -642
rect 1178 -643 1191 -638
rect 1178 -650 1182 -643
rect 1051 -660 1063 -650
rect 1095 -660 1106 -650
rect 1139 -660 1150 -650
rect 1039 -665 1043 -660
rect 1075 -665 1079 -660
rect 1119 -665 1123 -660
rect 1170 -665 1174 -660
rect 1038 -669 1182 -665
rect 802 -689 805 -683
rect 811 -711 814 -701
rect 791 -715 803 -711
rect 811 -714 823 -711
rect 895 -713 923 -710
rect 811 -719 814 -714
rect 896 -719 899 -713
rect 920 -714 923 -713
rect 920 -717 991 -714
rect 802 -743 805 -726
rect 879 -743 882 -740
rect 791 -746 805 -743
rect 887 -742 897 -739
rect 905 -739 908 -731
rect 935 -723 938 -717
rect 954 -723 957 -717
rect 905 -742 926 -739
rect 905 -745 908 -742
rect 896 -755 899 -751
rect 890 -757 914 -755
rect 890 -758 908 -757
rect 913 -758 914 -757
rect 923 -765 926 -742
rect 964 -723 984 -720
rect 964 -729 967 -723
rect 981 -729 984 -723
rect 945 -750 948 -747
rect 945 -753 963 -750
rect 1050 -739 1203 -735
rect 1056 -745 1060 -739
rect 1094 -745 1098 -739
rect 1138 -745 1142 -739
rect 1183 -745 1187 -739
rect 973 -760 976 -753
rect 973 -763 990 -760
rect 895 -766 914 -765
rect 890 -768 914 -766
rect 923 -768 966 -765
rect 896 -774 899 -768
rect 987 -774 990 -763
rect 1106 -770 1119 -745
rect 1150 -770 1163 -745
rect 952 -779 977 -776
rect 987 -778 1000 -774
rect 952 -781 955 -779
rect 794 -794 826 -791
rect 805 -800 808 -794
rect 879 -797 882 -794
rect 887 -797 897 -794
rect 905 -794 908 -786
rect 917 -784 955 -781
rect 987 -782 990 -778
rect 917 -794 920 -784
rect 958 -785 990 -782
rect 958 -788 961 -785
rect 905 -797 920 -794
rect 905 -800 908 -797
rect 957 -791 963 -788
rect 896 -810 899 -806
rect 917 -807 922 -804
rect 935 -804 938 -800
rect 982 -804 985 -800
rect 927 -807 991 -804
rect 917 -810 920 -807
rect 814 -822 817 -812
rect 890 -813 920 -810
rect 996 -818 1000 -778
rect 1045 -781 1052 -777
rect 1056 -789 1065 -785
rect 1072 -792 1076 -770
rect 1080 -781 1081 -777
rect 1116 -779 1119 -770
rect 1160 -779 1163 -770
rect 1116 -784 1128 -779
rect 1160 -784 1184 -779
rect 1191 -780 1195 -770
rect 1080 -786 1088 -784
rect 1085 -789 1088 -786
rect 1107 -789 1108 -785
rect 1116 -792 1119 -784
rect 1124 -789 1132 -784
rect 1151 -789 1152 -785
rect 1160 -792 1163 -784
rect 1191 -785 1204 -780
rect 1191 -792 1195 -785
rect 1064 -802 1076 -792
rect 1108 -802 1119 -792
rect 1152 -802 1163 -792
rect 1052 -807 1056 -802
rect 1088 -807 1092 -802
rect 1132 -807 1136 -802
rect 1183 -807 1187 -802
rect 1051 -811 1195 -807
rect 794 -826 806 -822
rect 814 -825 826 -822
rect 814 -830 817 -825
rect 666 -848 670 -846
rect 643 -853 670 -848
rect 700 -850 704 -845
rect 721 -850 725 -845
rect 738 -850 742 -845
rect 756 -850 760 -844
rect 700 -853 760 -850
rect 805 -854 808 -837
rect 904 -847 932 -844
rect 543 -860 561 -856
rect 794 -857 808 -854
rect 905 -853 908 -847
rect 929 -848 932 -847
rect 929 -851 1000 -848
rect 264 -869 417 -865
rect 795 -866 827 -863
rect 270 -875 274 -869
rect 308 -875 312 -869
rect 352 -875 356 -869
rect 397 -875 401 -869
rect 806 -872 809 -866
rect 320 -900 333 -875
rect 364 -900 377 -875
rect 888 -877 891 -874
rect 896 -876 906 -873
rect 914 -873 917 -865
rect 944 -857 947 -851
rect 963 -857 966 -851
rect 914 -876 935 -873
rect 914 -879 917 -876
rect 815 -894 818 -884
rect 905 -889 908 -885
rect 899 -891 923 -889
rect 899 -892 917 -891
rect 795 -898 807 -894
rect 815 -897 827 -894
rect 259 -911 266 -907
rect 270 -919 279 -915
rect 286 -922 290 -900
rect 294 -911 295 -907
rect 330 -909 333 -900
rect 374 -909 377 -900
rect 330 -914 342 -909
rect 374 -914 398 -909
rect 405 -910 409 -900
rect 815 -902 818 -897
rect 922 -892 923 -891
rect 932 -899 935 -876
rect 973 -857 993 -854
rect 973 -863 976 -857
rect 990 -863 993 -857
rect 1060 -862 1213 -858
rect 954 -884 957 -881
rect 954 -887 972 -884
rect 1066 -868 1070 -862
rect 1104 -868 1108 -862
rect 1148 -868 1152 -862
rect 1193 -868 1197 -862
rect 982 -894 985 -887
rect 1116 -893 1129 -868
rect 1160 -893 1173 -868
rect 982 -897 999 -894
rect 904 -900 923 -899
rect 899 -902 923 -900
rect 932 -902 975 -899
rect 905 -908 908 -902
rect 996 -908 999 -897
rect 1055 -904 1062 -900
rect 294 -916 302 -914
rect 299 -919 302 -916
rect 321 -919 322 -915
rect 330 -922 333 -914
rect 338 -919 346 -914
rect 365 -919 366 -915
rect 374 -922 377 -914
rect 405 -915 418 -910
rect 405 -922 409 -915
rect 278 -932 290 -922
rect 322 -932 333 -922
rect 366 -932 377 -922
rect 806 -926 809 -909
rect 961 -913 986 -910
rect 996 -912 1009 -908
rect 1066 -912 1075 -908
rect 961 -915 964 -913
rect 795 -929 809 -926
rect 888 -931 891 -928
rect 896 -931 906 -928
rect 914 -928 917 -920
rect 926 -918 964 -915
rect 996 -916 999 -912
rect 926 -928 929 -918
rect 967 -919 999 -916
rect 967 -922 970 -919
rect 914 -931 929 -928
rect 266 -937 270 -932
rect 302 -937 306 -932
rect 346 -937 350 -932
rect 397 -937 401 -932
rect 914 -934 917 -931
rect 265 -941 409 -937
rect 629 -938 782 -934
rect 635 -944 639 -938
rect 673 -944 677 -938
rect 717 -944 721 -938
rect 762 -944 766 -938
rect 966 -925 972 -922
rect 905 -944 908 -940
rect 926 -941 931 -938
rect 944 -938 947 -934
rect 991 -938 994 -934
rect 936 -941 1000 -938
rect 926 -944 929 -941
rect 685 -969 698 -944
rect 729 -969 742 -944
rect 899 -947 929 -944
rect 1005 -952 1009 -912
rect 1082 -915 1086 -893
rect 1090 -904 1091 -900
rect 1126 -902 1129 -893
rect 1170 -902 1173 -893
rect 1126 -907 1138 -902
rect 1170 -907 1194 -902
rect 1201 -903 1205 -893
rect 1090 -909 1098 -907
rect 1095 -912 1098 -909
rect 1117 -912 1118 -908
rect 1126 -915 1129 -907
rect 1134 -912 1142 -907
rect 1161 -912 1162 -908
rect 1170 -915 1173 -907
rect 1201 -908 1214 -903
rect 1201 -915 1205 -908
rect 1074 -925 1086 -915
rect 1118 -925 1129 -915
rect 1162 -925 1173 -915
rect 1062 -930 1066 -925
rect 1098 -930 1102 -925
rect 1142 -930 1146 -925
rect 1193 -930 1197 -925
rect 1061 -934 1205 -930
rect 624 -980 631 -976
rect 635 -988 644 -984
rect 651 -991 655 -969
rect 659 -980 660 -976
rect 695 -978 698 -969
rect 739 -978 742 -969
rect 695 -983 707 -978
rect 739 -983 763 -978
rect 770 -979 774 -969
rect 659 -985 667 -983
rect 664 -988 667 -985
rect 686 -988 687 -984
rect 695 -991 698 -983
rect 703 -988 711 -983
rect 730 -988 731 -984
rect 739 -991 742 -983
rect 770 -984 783 -979
rect 770 -991 774 -984
rect 643 -1001 655 -991
rect 687 -1001 698 -991
rect 731 -1001 742 -991
rect 909 -996 937 -993
rect 631 -1006 635 -1001
rect 667 -1006 671 -1001
rect 711 -1006 715 -1001
rect 762 -1006 766 -1001
rect 910 -1002 913 -996
rect 934 -997 937 -996
rect 934 -1000 1005 -997
rect 630 -1010 774 -1006
rect 893 -1026 896 -1023
rect 901 -1025 911 -1022
rect 919 -1022 922 -1014
rect 949 -1006 952 -1000
rect 968 -1006 971 -1000
rect 919 -1025 940 -1022
rect 919 -1028 922 -1025
rect 910 -1038 913 -1034
rect 904 -1040 928 -1038
rect 904 -1041 922 -1040
rect 927 -1041 928 -1040
rect 937 -1048 940 -1025
rect 978 -1006 998 -1003
rect 978 -1012 981 -1006
rect 995 -1012 998 -1006
rect 1065 -1009 1218 -1005
rect 959 -1033 962 -1030
rect 959 -1036 977 -1033
rect 1071 -1015 1075 -1009
rect 1109 -1015 1113 -1009
rect 1153 -1015 1157 -1009
rect 1198 -1015 1202 -1009
rect 987 -1043 990 -1036
rect 1121 -1040 1134 -1015
rect 1165 -1040 1178 -1015
rect 987 -1046 1004 -1043
rect 909 -1049 928 -1048
rect 904 -1051 928 -1049
rect 937 -1051 980 -1048
rect 910 -1057 913 -1051
rect 1001 -1057 1004 -1046
rect 1060 -1051 1067 -1047
rect 966 -1062 991 -1059
rect 1001 -1061 1014 -1057
rect 1071 -1059 1080 -1055
rect 966 -1064 969 -1062
rect 893 -1080 896 -1077
rect 901 -1080 911 -1077
rect 919 -1077 922 -1069
rect 931 -1067 969 -1064
rect 1001 -1065 1004 -1061
rect 931 -1077 934 -1067
rect 972 -1068 1004 -1065
rect 972 -1071 975 -1068
rect 919 -1080 934 -1077
rect 919 -1083 922 -1080
rect 971 -1074 977 -1071
rect 910 -1093 913 -1089
rect 931 -1090 936 -1087
rect 949 -1087 952 -1083
rect 996 -1087 999 -1083
rect 941 -1090 1005 -1087
rect 931 -1093 934 -1090
rect 904 -1096 934 -1093
rect 1010 -1101 1014 -1061
rect 1087 -1062 1091 -1040
rect 1095 -1051 1096 -1047
rect 1131 -1049 1134 -1040
rect 1175 -1049 1178 -1040
rect 1131 -1054 1143 -1049
rect 1175 -1054 1199 -1049
rect 1206 -1050 1210 -1040
rect 1095 -1056 1103 -1054
rect 1100 -1059 1103 -1056
rect 1122 -1059 1123 -1055
rect 1131 -1062 1134 -1054
rect 1139 -1059 1147 -1054
rect 1166 -1059 1167 -1055
rect 1175 -1062 1178 -1054
rect 1206 -1055 1219 -1050
rect 1206 -1062 1210 -1055
rect 1079 -1072 1091 -1062
rect 1123 -1072 1134 -1062
rect 1167 -1072 1178 -1062
rect 1067 -1077 1071 -1072
rect 1103 -1077 1107 -1072
rect 1147 -1077 1151 -1072
rect 1198 -1077 1202 -1072
rect 1066 -1081 1210 -1077
<< m2contact >>
rect 509 -481 514 -476
rect 649 -481 654 -476
rect 66 -530 71 -525
rect 96 -522 101 -517
rect 95 -532 100 -527
rect 123 -530 128 -525
rect 167 -530 172 -525
rect 261 -527 266 -522
rect 291 -519 296 -514
rect 784 -481 789 -476
rect 922 -482 927 -477
rect 290 -529 295 -524
rect 318 -527 323 -522
rect 362 -527 367 -522
rect 509 -535 514 -530
rect 649 -535 654 -530
rect 784 -535 789 -530
rect 922 -536 927 -531
rect 63 -631 68 -626
rect 93 -623 98 -618
rect 92 -633 97 -628
rect 120 -631 125 -626
rect 164 -631 169 -626
rect 263 -625 268 -620
rect 293 -617 298 -612
rect 292 -627 297 -622
rect 320 -625 325 -620
rect 364 -625 369 -620
rect 871 -608 876 -603
rect 62 -728 67 -723
rect 92 -720 97 -715
rect 91 -730 96 -725
rect 119 -728 124 -723
rect 163 -728 168 -723
rect 262 -722 267 -717
rect 292 -714 297 -709
rect 291 -724 296 -719
rect 319 -722 324 -717
rect 363 -722 368 -717
rect 63 -824 68 -819
rect 93 -816 98 -811
rect 92 -826 97 -821
rect 120 -824 125 -819
rect 164 -824 169 -819
rect 263 -818 268 -813
rect 293 -810 298 -805
rect 292 -820 297 -815
rect 320 -818 325 -813
rect 364 -818 369 -813
rect 871 -662 876 -657
rect 1038 -647 1043 -642
rect 1068 -639 1073 -634
rect 1067 -649 1072 -644
rect 1095 -647 1100 -642
rect 1139 -647 1144 -642
rect 882 -744 887 -739
rect 882 -798 887 -793
rect 1051 -789 1056 -784
rect 1081 -781 1086 -776
rect 1080 -791 1085 -786
rect 1108 -789 1113 -784
rect 1152 -789 1157 -784
rect 891 -878 896 -873
rect 265 -919 270 -914
rect 295 -911 300 -906
rect 294 -921 299 -916
rect 322 -919 327 -914
rect 366 -919 371 -914
rect 1061 -912 1066 -907
rect 891 -932 896 -927
rect 1091 -904 1096 -899
rect 1090 -914 1095 -909
rect 1118 -912 1123 -907
rect 1162 -912 1167 -907
rect 630 -988 635 -983
rect 660 -980 665 -975
rect 659 -990 664 -985
rect 687 -988 692 -983
rect 731 -988 736 -983
rect 896 -1027 901 -1022
rect 1066 -1059 1071 -1054
rect 896 -1081 901 -1076
rect 1096 -1051 1101 -1046
rect 1095 -1061 1100 -1056
rect 1123 -1059 1128 -1054
rect 1167 -1059 1172 -1054
<< pm12contact >>
rect 565 -498 570 -493
rect 574 -499 579 -494
rect 705 -498 710 -493
rect 714 -499 719 -494
rect 840 -498 845 -493
rect 849 -499 854 -494
rect 978 -499 983 -494
rect 987 -500 992 -495
rect 927 -625 932 -620
rect 936 -626 941 -621
rect 938 -761 943 -756
rect 947 -762 952 -757
rect 947 -895 952 -890
rect 956 -896 961 -891
rect 952 -1044 957 -1039
rect 961 -1045 966 -1040
<< metal2 >>
rect 291 -469 322 -466
rect 96 -472 127 -469
rect 96 -517 100 -472
rect 123 -525 127 -472
rect 291 -514 295 -469
rect 318 -522 322 -469
rect 510 -487 513 -481
rect 650 -487 653 -481
rect 785 -487 788 -481
rect 510 -490 547 -487
rect 650 -490 687 -487
rect 785 -490 822 -487
rect 544 -493 547 -490
rect 684 -493 687 -490
rect 819 -493 822 -490
rect 923 -488 926 -482
rect 923 -491 960 -488
rect 544 -496 565 -493
rect 574 -509 577 -499
rect 684 -496 705 -493
rect 714 -509 717 -499
rect 819 -496 840 -493
rect 957 -494 960 -491
rect 849 -509 852 -499
rect 957 -497 978 -494
rect 511 -512 577 -509
rect 651 -512 717 -509
rect 786 -512 852 -509
rect 987 -510 990 -500
rect 45 -530 66 -526
rect 57 -554 63 -530
rect 240 -527 261 -523
rect 96 -554 100 -532
rect 167 -554 172 -530
rect 252 -551 258 -527
rect 291 -551 295 -529
rect 362 -551 367 -527
rect 511 -530 514 -512
rect 651 -530 654 -512
rect 786 -530 789 -512
rect 924 -513 990 -510
rect 924 -531 927 -513
rect 252 -554 371 -551
rect 57 -557 176 -554
rect 293 -567 324 -564
rect 93 -573 124 -570
rect 93 -618 97 -573
rect 120 -626 124 -573
rect 293 -612 297 -567
rect 320 -620 324 -567
rect 1068 -589 1099 -586
rect 872 -614 875 -608
rect 872 -617 909 -614
rect 906 -620 909 -617
rect 242 -625 263 -621
rect 42 -631 63 -627
rect 54 -655 60 -631
rect 93 -655 97 -633
rect 164 -655 169 -631
rect 254 -649 260 -625
rect 293 -649 297 -627
rect 364 -649 369 -625
rect 906 -623 927 -620
rect 936 -636 939 -626
rect 873 -639 939 -636
rect 1068 -634 1072 -589
rect 254 -652 373 -649
rect 54 -658 173 -655
rect 873 -657 876 -639
rect 1095 -642 1099 -589
rect 1017 -647 1038 -643
rect 292 -664 323 -661
rect 92 -670 123 -667
rect 92 -715 96 -670
rect 119 -723 123 -670
rect 292 -709 296 -664
rect 319 -717 323 -664
rect 1029 -671 1035 -647
rect 1068 -671 1072 -649
rect 1139 -671 1144 -647
rect 1029 -674 1148 -671
rect 241 -722 262 -718
rect 41 -728 62 -724
rect 53 -752 59 -728
rect 92 -752 96 -730
rect 163 -752 168 -728
rect 253 -746 259 -722
rect 292 -746 296 -724
rect 363 -746 368 -722
rect 1081 -731 1112 -728
rect 253 -749 372 -746
rect 883 -750 886 -744
rect 53 -755 172 -752
rect 883 -753 920 -750
rect 917 -756 920 -753
rect 293 -760 324 -757
rect 93 -766 124 -763
rect 93 -811 97 -766
rect 120 -819 124 -766
rect 293 -805 297 -760
rect 320 -813 324 -760
rect 917 -759 938 -756
rect 947 -772 950 -762
rect 884 -775 950 -772
rect 884 -793 887 -775
rect 1081 -776 1085 -731
rect 1108 -784 1112 -731
rect 1030 -789 1051 -785
rect 1042 -813 1048 -789
rect 1081 -813 1085 -791
rect 1152 -813 1157 -789
rect 242 -818 263 -814
rect 42 -824 63 -820
rect 54 -848 60 -824
rect 93 -848 97 -826
rect 164 -848 169 -824
rect 254 -842 260 -818
rect 1042 -816 1161 -813
rect 293 -842 297 -820
rect 364 -842 369 -818
rect 254 -845 373 -842
rect 54 -851 173 -848
rect 1091 -854 1122 -851
rect 295 -861 326 -858
rect 295 -906 299 -861
rect 322 -914 326 -861
rect 892 -884 895 -878
rect 892 -887 929 -884
rect 926 -890 929 -887
rect 926 -893 947 -890
rect 956 -906 959 -896
rect 1091 -899 1095 -854
rect 893 -909 959 -906
rect 1118 -907 1122 -854
rect 244 -919 265 -915
rect 256 -943 262 -919
rect 295 -943 299 -921
rect 366 -943 371 -919
rect 893 -927 896 -909
rect 1040 -912 1061 -908
rect 660 -930 691 -927
rect 256 -946 375 -943
rect 660 -975 664 -930
rect 687 -983 691 -930
rect 1052 -936 1058 -912
rect 1091 -936 1095 -914
rect 1162 -936 1167 -912
rect 1052 -939 1171 -936
rect 609 -988 630 -984
rect 621 -1012 627 -988
rect 660 -1012 664 -990
rect 731 -1012 736 -988
rect 1096 -1001 1127 -998
rect 621 -1015 740 -1012
rect 897 -1033 900 -1027
rect 897 -1036 934 -1033
rect 931 -1039 934 -1036
rect 931 -1042 952 -1039
rect 961 -1055 964 -1045
rect 1096 -1046 1100 -1001
rect 1123 -1054 1127 -1001
rect 898 -1058 964 -1055
rect 898 -1076 901 -1058
rect 1045 -1059 1066 -1055
rect 1057 -1083 1063 -1059
rect 1096 -1083 1100 -1061
rect 1167 -1083 1172 -1059
rect 1057 -1086 1176 -1083
<< m123contact >>
rect 517 -450 522 -445
rect 657 -450 662 -445
rect 792 -450 797 -445
rect 930 -451 935 -446
rect 517 -503 522 -498
rect 535 -499 540 -494
rect 657 -503 662 -498
rect 675 -499 680 -494
rect 792 -503 797 -498
rect 810 -499 815 -494
rect 930 -504 935 -499
rect 948 -500 953 -495
rect 549 -544 554 -539
rect 689 -544 694 -539
rect 824 -544 829 -539
rect 962 -545 967 -540
rect 879 -577 884 -572
rect 879 -630 884 -625
rect 897 -626 902 -621
rect 911 -671 916 -666
rect 890 -713 895 -708
rect 890 -766 895 -761
rect 908 -762 913 -757
rect 922 -807 927 -802
rect 899 -847 904 -842
rect 899 -900 904 -895
rect 917 -896 922 -891
rect 931 -941 936 -936
rect 904 -996 909 -991
rect 904 -1049 909 -1044
rect 922 -1045 927 -1040
rect 936 -1090 941 -1085
<< metal3 >>
rect 517 -498 520 -450
rect 540 -499 552 -496
rect 549 -539 552 -499
rect 657 -498 660 -450
rect 680 -499 692 -496
rect 689 -539 692 -499
rect 792 -498 795 -450
rect 815 -499 827 -496
rect 824 -539 827 -499
rect 930 -499 933 -451
rect 953 -500 965 -497
rect 962 -540 965 -500
rect 879 -625 882 -577
rect 902 -626 914 -623
rect 911 -666 914 -626
rect 890 -761 893 -713
rect 913 -762 925 -759
rect 922 -802 925 -762
rect 899 -895 902 -847
rect 922 -896 934 -893
rect 931 -936 934 -896
rect 904 -1044 907 -996
rect 927 -1045 939 -1042
rect 936 -1085 939 -1045
<< labels >>
rlabel metal1 535 -550 539 -547 1 gnd
rlabel metal1 585 -544 588 -542 1 gnd
rlabel metal1 533 -494 534 -492 1 gnd
rlabel metal1 529 -450 532 -448 5 vdd
rlabel metal1 530 -504 533 -502 1 vdd
rlabel metal1 614 -515 618 -511 7 p0
rlabel metal1 506 -480 507 -477 1 a0
rlabel metal1 506 -534 507 -531 1 b0
rlabel metal1 675 -550 679 -547 1 gnd
rlabel metal1 725 -544 728 -542 1 gnd
rlabel metal1 673 -494 674 -492 1 gnd
rlabel metal1 669 -450 672 -448 5 vdd
rlabel metal1 670 -504 673 -502 1 vdd
rlabel metal1 810 -550 814 -547 1 gnd
rlabel metal1 860 -544 863 -542 1 gnd
rlabel metal1 808 -494 809 -492 1 gnd
rlabel metal1 804 -450 807 -448 5 vdd
rlabel metal1 805 -504 808 -502 1 vdd
rlabel metal1 948 -551 952 -548 1 gnd
rlabel metal1 998 -545 1001 -543 1 gnd
rlabel metal1 946 -495 947 -493 1 gnd
rlabel metal1 942 -451 945 -449 5 vdd
rlabel metal1 943 -505 946 -503 1 vdd
rlabel metal1 646 -534 647 -531 1 b1
rlabel metal1 646 -480 647 -477 1 a1
rlabel metal1 781 -480 782 -477 1 a2
rlabel metal1 781 -534 782 -531 1 b2
rlabel metal1 919 -481 920 -478 1 a3
rlabel metal1 919 -535 920 -532 1 b3
rlabel metal1 1027 -516 1031 -512 7 p3
rlabel metal1 754 -515 758 -511 1 p1
rlabel metal1 889 -515 893 -511 1 p2
rlabel metal1 508 -605 509 -604 7 g0
rlabel metal1 445 -611 446 -610 3 b0
rlabel metal1 443 -604 444 -603 3 a0
rlabel metal1 468 -637 468 -637 1 gnd!
rlabel metal1 468 -573 468 -573 5 vdd!
rlabel metal1 508 -679 509 -678 7 g1
rlabel metal1 468 -780 468 -780 1 gnd!
rlabel metal1 468 -716 468 -716 5 vdd!
rlabel metal1 468 -854 468 -854 1 gnd!
rlabel metal1 468 -790 468 -790 5 vdd!
rlabel metal1 443 -747 444 -746 3 a2
rlabel metal1 445 -754 446 -753 3 b2
rlabel metal1 444 -821 445 -820 3 a3
rlabel metal1 445 -828 446 -827 3 b3
rlabel metal1 508 -822 509 -821 7 g3
rlabel metal1 445 -685 446 -684 3 b1
rlabel metal1 444 -678 445 -677 3 a1
rlabel metal1 468 -647 468 -647 5 vdd!
rlabel metal1 468 -711 468 -711 1 gnd!
rlabel metal1 561 -572 568 -571 1 vdd
rlabel metal1 550 -605 553 -603 1 gnd
rlabel metal1 565 -604 566 -603 1 c3b
rlabel metal1 547 -618 548 -617 1 cin
rlabel metal1 568 -618 569 -616 1 p0
rlabel metal1 597 -572 604 -571 1 vdd
rlabel metal1 586 -605 589 -603 1 gnd
rlabel metal1 638 -572 645 -571 1 vdd
rlabel metal1 627 -605 630 -603 1 gnd
rlabel metal1 673 -572 680 -571 1 vdd
rlabel metal1 662 -605 665 -603 1 gnd
rlabel metal1 601 -604 602 -603 1 c2b
rlabel metal1 642 -604 643 -603 1 c1b
rlabel metal1 677 -604 678 -603 1 c0b
rlabel metal1 601 -618 602 -617 1 p1
rlabel metal1 634 -618 635 -617 1 p2
rlabel metal1 665 -618 666 -617 1 p3
rlabel metal1 675 -619 677 -617 1 c3b
rlabel metal1 699 -617 700 -616 1 g0
rlabel metal1 709 -618 711 -616 1 c0b
rlabel metal1 720 -617 721 -616 1 g1
rlabel metal1 730 -618 732 -616 1 c1b
rlabel metal1 737 -617 738 -616 1 g2
rlabel metal1 747 -618 749 -616 1 c2b
rlabel metal1 755 -616 756 -615 1 g3
rlabel metal1 765 -617 767 -615 1 c3b
rlabel metal1 897 -677 901 -674 1 gnd
rlabel metal1 947 -671 950 -669 1 gnd
rlabel metal1 895 -621 896 -619 1 gnd
rlabel metal1 891 -577 894 -575 5 vdd
rlabel metal1 892 -631 895 -629 1 vdd
rlabel metal1 908 -813 912 -810 1 gnd
rlabel metal1 958 -807 961 -805 1 gnd
rlabel metal1 906 -757 907 -755 1 gnd
rlabel metal1 902 -713 905 -711 5 vdd
rlabel metal1 903 -767 906 -765 1 vdd
rlabel metal1 917 -947 921 -944 1 gnd
rlabel metal1 967 -941 970 -939 1 gnd
rlabel metal1 915 -891 916 -889 1 gnd
rlabel metal1 911 -847 914 -845 5 vdd
rlabel metal1 912 -901 915 -899 1 vdd
rlabel metal1 922 -1096 926 -1093 1 gnd
rlabel metal1 972 -1090 975 -1088 1 gnd
rlabel metal1 920 -1040 921 -1038 1 gnd
rlabel metal1 916 -996 919 -994 5 vdd
rlabel metal1 917 -1050 920 -1048 1 vdd
rlabel metal1 868 -607 869 -604 1 p0
rlabel metal1 868 -661 869 -658 1 cin
rlabel metal1 976 -642 980 -638 1 s0
rlabel metal1 879 -743 880 -740 1 p1
rlabel metal1 879 -797 880 -794 1 c0
rlabel metal1 987 -778 991 -774 1 s1
rlabel metal1 888 -877 889 -874 1 p2
rlabel metal1 888 -931 889 -928 1 c1
rlabel metal1 996 -912 1000 -908 1 s2
rlabel metal1 893 -1026 894 -1023 1 p3
rlabel metal1 893 -1080 894 -1077 1 c2
rlabel metal1 1001 -1061 1005 -1057 1 s3
rlabel metal1 508 -748 509 -747 7 g2
rlabel metal1 793 -629 794 -627 1 c0b
rlabel metal1 795 -714 798 -712 1 c1b
rlabel metal1 799 -825 802 -823 1 c2b
rlabel metal1 800 -897 803 -895 1 c3b
rlabel metal1 817 -628 820 -626 1 c0
rlabel metal1 818 -713 819 -712 1 c1
rlabel metal1 821 -824 822 -823 1 c2
rlabel metal1 822 -896 823 -895 1 c3
rlabel metal1 800 -928 802 -927 1 gnd
rlabel metal1 807 -865 809 -864 1 vdd
rlabel metal1 800 -855 802 -854 1 gnd
rlabel metal1 806 -793 808 -792 1 vdd
rlabel metal1 797 -745 799 -744 1 gnd
rlabel metal1 805 -682 807 -681 1 vdd
rlabel metal1 794 -660 796 -659 1 gnd
rlabel metal1 802 -597 804 -596 1 vdd
rlabel metal1 270 -547 273 -546 1 gnd
rlabel metal1 276 -475 278 -474 5 vdd
rlabel metal2 259 -525 261 -524 1 clk
rlabel metal1 408 -523 411 -519 1 a0
rlabel metal1 257 -518 259 -516 1 a0d
rlabel metal1 272 -645 275 -644 1 gnd
rlabel metal1 278 -573 280 -572 5 vdd
rlabel metal2 261 -623 263 -622 1 clk
rlabel metal1 271 -742 274 -741 1 gnd
rlabel metal1 277 -670 279 -669 5 vdd
rlabel metal2 260 -720 262 -719 1 clk
rlabel metal1 272 -838 275 -837 1 gnd
rlabel metal1 278 -766 280 -765 5 vdd
rlabel metal2 261 -816 263 -815 1 clk
rlabel metal1 75 -550 78 -549 1 gnd
rlabel metal1 81 -478 83 -477 5 vdd
rlabel metal2 64 -528 66 -527 1 clk
rlabel metal2 61 -822 63 -821 1 clk
rlabel metal1 78 -772 80 -771 5 vdd
rlabel metal1 72 -844 75 -843 1 gnd
rlabel metal2 60 -726 62 -725 1 clk
rlabel metal1 77 -676 79 -675 5 vdd
rlabel metal1 71 -748 74 -747 1 gnd
rlabel metal2 61 -629 63 -628 1 clk
rlabel metal1 78 -579 80 -578 5 vdd
rlabel metal1 72 -651 75 -650 1 gnd
rlabel metal1 62 -521 64 -519 1 b0d
rlabel metal1 213 -526 216 -522 1 b0
rlabel metal1 59 -622 61 -620 1 b1d
rlabel metal1 210 -627 213 -623 1 b1
rlabel metal1 58 -719 60 -717 1 b2d
rlabel metal1 209 -724 212 -720 1 b2
rlabel metal1 59 -815 61 -813 1 b3d
rlabel metal1 210 -820 213 -816 1 b3
rlabel metal1 410 -621 413 -617 1 a1
rlabel metal1 259 -616 261 -614 1 a1d
rlabel metal1 258 -713 260 -711 1 a2d
rlabel metal1 409 -718 412 -714 1 a2
rlabel metal1 259 -809 261 -807 1 a3d
rlabel metal1 410 -814 413 -810 1 a3
rlabel metal1 274 -939 277 -938 1 gnd
rlabel metal1 280 -867 282 -866 5 vdd
rlabel metal2 263 -917 265 -916 1 clk
rlabel metal1 412 -915 415 -911 1 cin
rlabel metal1 261 -909 263 -908 1 cind
rlabel metal1 1047 -667 1050 -666 1 gnd
rlabel metal1 1053 -595 1055 -594 5 vdd
rlabel metal2 1036 -645 1038 -644 1 clk
rlabel metal1 1060 -809 1063 -808 1 gnd
rlabel metal1 1066 -737 1068 -736 5 vdd
rlabel metal2 1049 -787 1051 -786 1 clk
rlabel metal1 1070 -932 1073 -931 1 gnd
rlabel metal1 1076 -860 1078 -859 5 vdd
rlabel metal2 1059 -910 1061 -909 1 clk
rlabel metal1 1075 -1079 1078 -1078 1 gnd
rlabel metal1 1081 -1007 1083 -1006 5 vdd
rlabel metal2 1064 -1057 1066 -1056 1 clk
rlabel metal1 1062 -1050 1064 -1048 1 s3
rlabel metal1 1213 -1055 1216 -1051 7 s3d
rlabel metal1 1208 -908 1211 -904 1 s2d
rlabel metal1 1057 -903 1059 -901 1 s2
rlabel metal1 1047 -780 1049 -778 1 s1
rlabel metal1 1034 -638 1037 -636 1 s0
rlabel metal1 1184 -643 1189 -639 1 s0d
rlabel metal1 1198 -785 1201 -781 1 s1d
rlabel metal1 723 -853 726 -851 1 gnd
rlabel metal1 654 -853 661 -848 1 c2b
rlabel metal1 619 -853 626 -848 1 c1b
rlabel metal1 580 -853 587 -848 1 c0b
rlabel metal1 552 -859 558 -857 1 gnd
rlabel metal1 639 -1008 642 -1007 1 gnd
rlabel metal1 645 -936 647 -935 5 vdd
rlabel metal2 628 -986 630 -985 1 clk
rlabel metal1 626 -979 628 -977 1 c3
rlabel metal1 777 -984 780 -980 1 coutd
<< end >>
