magic
tech scmos
timestamp 1731729581
<< nwell >>
rect 177 180 201 204
rect 216 194 250 200
rect 216 164 278 194
rect 317 180 341 204
rect 356 194 390 200
rect 356 164 418 194
rect 452 180 476 204
rect 491 194 525 200
rect 491 164 553 194
rect 590 179 614 203
rect 629 193 663 199
rect 244 158 278 164
rect 384 158 418 164
rect 519 158 553 164
rect 629 163 691 193
rect 657 157 691 163
rect 177 125 201 149
rect 317 125 341 149
rect 452 125 476 149
rect 590 124 614 148
rect 102 53 139 79
rect 145 53 173 79
rect 208 55 236 81
rect 244 55 272 81
rect 285 55 313 81
rect 320 55 348 81
rect 454 30 482 56
rect 539 53 563 77
rect 578 67 612 73
rect 578 37 640 67
rect 606 31 640 37
rect 102 -21 139 5
rect 145 -21 173 5
rect 539 -2 563 22
rect 455 -55 483 -29
rect 102 -90 139 -64
rect 145 -90 173 -64
rect 550 -83 574 -59
rect 589 -69 623 -63
rect 589 -99 651 -69
rect 617 -105 651 -99
rect 550 -138 574 -114
rect 102 -164 139 -138
rect 145 -164 173 -138
rect 458 -166 486 -140
rect 459 -238 487 -212
rect 559 -217 583 -193
rect 598 -203 632 -197
rect 598 -233 660 -203
rect 626 -239 660 -233
rect 559 -272 583 -248
rect 564 -366 588 -342
rect 603 -352 637 -346
rect 603 -382 665 -352
rect 631 -388 665 -382
rect 564 -421 588 -397
<< ntransistor >>
rect 188 166 190 172
rect 328 166 330 172
rect 463 166 465 172
rect 227 117 229 129
rect 237 117 239 129
rect 255 117 257 129
rect 265 117 267 129
rect 601 165 603 171
rect 367 117 369 129
rect 377 117 379 129
rect 395 117 397 129
rect 405 117 407 129
rect 502 117 504 129
rect 512 117 514 129
rect 530 117 532 129
rect 540 117 542 129
rect 188 111 190 117
rect 328 111 330 117
rect 463 111 465 117
rect 640 116 642 128
rect 650 116 652 128
rect 668 116 670 128
rect 678 116 680 128
rect 601 110 603 116
rect 115 25 117 38
rect 125 25 127 38
rect 157 36 159 43
rect 550 39 552 45
rect 115 -49 117 -36
rect 125 -49 127 -36
rect 157 -38 159 -31
rect 115 -118 117 -105
rect 125 -118 127 -105
rect 157 -107 159 -100
rect 115 -192 117 -179
rect 125 -192 127 -179
rect 157 -181 159 -174
rect 213 -229 215 31
rect 220 -229 222 31
rect 267 -228 269 32
rect 300 -228 302 32
rect 331 -228 333 32
rect 365 -227 367 33
rect 386 -227 388 33
rect 403 -227 405 33
rect 421 -226 423 34
rect 466 13 468 20
rect 589 -10 591 2
rect 599 -10 601 2
rect 617 -10 619 2
rect 627 -10 629 2
rect 550 -16 552 -10
rect 467 -72 469 -65
rect 561 -97 563 -91
rect 600 -146 602 -134
rect 610 -146 612 -134
rect 628 -146 630 -134
rect 638 -146 640 -134
rect 561 -152 563 -146
rect 470 -183 472 -176
rect 570 -231 572 -225
rect 471 -255 473 -248
rect 609 -280 611 -268
rect 619 -280 621 -268
rect 637 -280 639 -268
rect 647 -280 649 -268
rect 570 -286 572 -280
rect 575 -380 577 -374
rect 614 -429 616 -417
rect 624 -429 626 -417
rect 642 -429 644 -417
rect 652 -429 654 -417
rect 575 -435 577 -429
<< ptransistor >>
rect 188 186 190 198
rect 227 170 229 194
rect 237 170 239 194
rect 255 164 257 188
rect 265 164 267 188
rect 328 186 330 198
rect 367 170 369 194
rect 377 170 379 194
rect 188 131 190 143
rect 395 164 397 188
rect 405 164 407 188
rect 463 186 465 198
rect 502 170 504 194
rect 512 170 514 194
rect 328 131 330 143
rect 530 164 532 188
rect 540 164 542 188
rect 601 185 603 197
rect 640 169 642 193
rect 650 169 652 193
rect 463 131 465 143
rect 668 163 670 187
rect 678 163 680 187
rect 601 130 603 142
rect 115 61 117 73
rect 125 61 127 73
rect 157 61 159 73
rect 220 63 222 75
rect 256 63 258 75
rect 297 63 299 75
rect 332 63 334 75
rect 550 59 552 71
rect 466 38 468 50
rect 589 43 591 67
rect 599 43 601 67
rect 115 -13 117 -1
rect 125 -13 127 -1
rect 157 -13 159 -1
rect 115 -82 117 -70
rect 125 -82 127 -70
rect 157 -82 159 -70
rect 115 -156 117 -144
rect 125 -156 127 -144
rect 157 -156 159 -144
rect 617 37 619 61
rect 627 37 629 61
rect 550 4 552 16
rect 467 -47 469 -35
rect 561 -77 563 -65
rect 600 -93 602 -69
rect 610 -93 612 -69
rect 628 -99 630 -75
rect 638 -99 640 -75
rect 561 -132 563 -120
rect 470 -158 472 -146
rect 570 -211 572 -199
rect 471 -230 473 -218
rect 609 -227 611 -203
rect 619 -227 621 -203
rect 637 -233 639 -209
rect 647 -233 649 -209
rect 570 -266 572 -254
rect 575 -360 577 -348
rect 614 -376 616 -352
rect 624 -376 626 -352
rect 642 -382 644 -358
rect 652 -382 654 -358
rect 575 -415 577 -403
<< ndiffusion >>
rect 187 166 188 172
rect 190 166 191 172
rect 327 166 328 172
rect 330 166 331 172
rect 462 166 463 172
rect 465 166 466 172
rect 226 117 227 129
rect 229 117 237 129
rect 239 117 240 129
rect 254 117 255 129
rect 257 117 265 129
rect 267 117 268 129
rect 600 165 601 171
rect 603 165 604 171
rect 366 117 367 129
rect 369 117 377 129
rect 379 117 380 129
rect 394 117 395 129
rect 397 117 405 129
rect 407 117 408 129
rect 501 117 502 129
rect 504 117 512 129
rect 514 117 515 129
rect 529 117 530 129
rect 532 117 540 129
rect 542 117 543 129
rect 187 111 188 117
rect 190 111 191 117
rect 327 111 328 117
rect 330 111 331 117
rect 462 111 463 117
rect 465 111 466 117
rect 639 116 640 128
rect 642 116 650 128
rect 652 116 653 128
rect 667 116 668 128
rect 670 116 678 128
rect 680 116 681 128
rect 600 110 601 116
rect 603 110 604 116
rect 114 25 115 38
rect 117 25 125 38
rect 127 25 128 38
rect 156 36 157 43
rect 159 36 160 43
rect 549 39 550 45
rect 552 39 553 45
rect 114 -49 115 -36
rect 117 -49 125 -36
rect 127 -49 128 -36
rect 156 -38 157 -31
rect 159 -38 160 -31
rect 114 -118 115 -105
rect 117 -118 125 -105
rect 127 -118 128 -105
rect 156 -107 157 -100
rect 159 -107 160 -100
rect 114 -192 115 -179
rect 117 -192 125 -179
rect 127 -192 128 -179
rect 156 -181 157 -174
rect 159 -181 160 -174
rect 212 -229 213 31
rect 215 -229 220 31
rect 222 -229 223 31
rect 266 -228 267 32
rect 269 -228 270 32
rect 299 -228 300 32
rect 302 -228 303 32
rect 330 -228 331 32
rect 333 -228 334 32
rect 364 -227 365 33
rect 367 -227 368 33
rect 385 -227 386 33
rect 388 -227 389 33
rect 402 -227 403 33
rect 405 -227 406 33
rect 420 -226 421 34
rect 423 -226 424 34
rect 465 13 466 20
rect 468 13 469 20
rect 588 -10 589 2
rect 591 -10 599 2
rect 601 -10 602 2
rect 616 -10 617 2
rect 619 -10 627 2
rect 629 -10 630 2
rect 549 -16 550 -10
rect 552 -16 553 -10
rect 466 -72 467 -65
rect 469 -72 470 -65
rect 560 -97 561 -91
rect 563 -97 564 -91
rect 599 -146 600 -134
rect 602 -146 610 -134
rect 612 -146 613 -134
rect 627 -146 628 -134
rect 630 -146 638 -134
rect 640 -146 641 -134
rect 560 -152 561 -146
rect 563 -152 564 -146
rect 469 -183 470 -176
rect 472 -183 473 -176
rect 569 -231 570 -225
rect 572 -231 573 -225
rect 470 -255 471 -248
rect 473 -255 474 -248
rect 608 -280 609 -268
rect 611 -280 619 -268
rect 621 -280 622 -268
rect 636 -280 637 -268
rect 639 -280 647 -268
rect 649 -280 650 -268
rect 569 -286 570 -280
rect 572 -286 573 -280
rect 574 -380 575 -374
rect 577 -380 578 -374
rect 613 -429 614 -417
rect 616 -429 624 -417
rect 626 -429 627 -417
rect 641 -429 642 -417
rect 644 -429 652 -417
rect 654 -429 655 -417
rect 574 -435 575 -429
rect 577 -435 578 -429
<< pdiffusion >>
rect 187 186 188 198
rect 190 186 191 198
rect 226 170 227 194
rect 229 170 231 194
rect 235 170 237 194
rect 239 170 240 194
rect 254 164 255 188
rect 257 164 259 188
rect 263 164 265 188
rect 267 164 268 188
rect 327 186 328 198
rect 330 186 331 198
rect 366 170 367 194
rect 369 170 371 194
rect 375 170 377 194
rect 379 170 380 194
rect 187 131 188 143
rect 190 131 191 143
rect 394 164 395 188
rect 397 164 399 188
rect 403 164 405 188
rect 407 164 408 188
rect 462 186 463 198
rect 465 186 466 198
rect 501 170 502 194
rect 504 170 506 194
rect 510 170 512 194
rect 514 170 515 194
rect 327 131 328 143
rect 330 131 331 143
rect 529 164 530 188
rect 532 164 534 188
rect 538 164 540 188
rect 542 164 543 188
rect 600 185 601 197
rect 603 185 604 197
rect 639 169 640 193
rect 642 169 644 193
rect 648 169 650 193
rect 652 169 653 193
rect 462 131 463 143
rect 465 131 466 143
rect 667 163 668 187
rect 670 163 672 187
rect 676 163 678 187
rect 680 163 681 187
rect 600 130 601 142
rect 603 130 604 142
rect 114 61 115 73
rect 117 61 119 73
rect 123 61 125 73
rect 127 61 128 73
rect 156 61 157 73
rect 159 61 160 73
rect 219 63 220 75
rect 222 63 223 75
rect 255 63 256 75
rect 258 63 259 75
rect 296 63 297 75
rect 299 63 300 75
rect 331 63 332 75
rect 334 63 335 75
rect 549 59 550 71
rect 552 59 553 71
rect 465 38 466 50
rect 468 38 469 50
rect 588 43 589 67
rect 591 43 593 67
rect 597 43 599 67
rect 601 43 602 67
rect 114 -13 115 -1
rect 117 -13 119 -1
rect 123 -13 125 -1
rect 127 -13 128 -1
rect 156 -13 157 -1
rect 159 -13 160 -1
rect 114 -82 115 -70
rect 117 -82 119 -70
rect 123 -82 125 -70
rect 127 -82 128 -70
rect 156 -82 157 -70
rect 159 -82 160 -70
rect 114 -156 115 -144
rect 117 -156 119 -144
rect 123 -156 125 -144
rect 127 -156 128 -144
rect 156 -156 157 -144
rect 159 -156 160 -144
rect 616 37 617 61
rect 619 37 621 61
rect 625 37 627 61
rect 629 37 630 61
rect 549 4 550 16
rect 552 4 553 16
rect 466 -47 467 -35
rect 469 -47 470 -35
rect 560 -77 561 -65
rect 563 -77 564 -65
rect 599 -93 600 -69
rect 602 -93 604 -69
rect 608 -93 610 -69
rect 612 -93 613 -69
rect 627 -99 628 -75
rect 630 -99 632 -75
rect 636 -99 638 -75
rect 640 -99 641 -75
rect 560 -132 561 -120
rect 563 -132 564 -120
rect 469 -158 470 -146
rect 472 -158 473 -146
rect 569 -211 570 -199
rect 572 -211 573 -199
rect 470 -230 471 -218
rect 473 -230 474 -218
rect 608 -227 609 -203
rect 611 -227 613 -203
rect 617 -227 619 -203
rect 621 -227 622 -203
rect 636 -233 637 -209
rect 639 -233 641 -209
rect 645 -233 647 -209
rect 649 -233 650 -209
rect 569 -266 570 -254
rect 572 -266 573 -254
rect 574 -360 575 -348
rect 577 -360 578 -348
rect 613 -376 614 -352
rect 616 -376 618 -352
rect 622 -376 624 -352
rect 626 -376 627 -352
rect 641 -382 642 -358
rect 644 -382 646 -358
rect 650 -382 652 -358
rect 654 -382 655 -358
rect 574 -415 575 -403
rect 577 -415 578 -403
<< ndcontact >>
rect 183 166 187 172
rect 191 166 195 172
rect 323 166 327 172
rect 331 166 335 172
rect 458 166 462 172
rect 466 166 470 172
rect 222 117 226 129
rect 240 117 244 129
rect 250 117 254 129
rect 268 117 272 129
rect 596 165 600 171
rect 604 165 608 171
rect 362 117 366 129
rect 380 117 384 129
rect 390 117 394 129
rect 408 117 412 129
rect 497 117 501 129
rect 515 117 519 129
rect 525 117 529 129
rect 543 117 547 129
rect 183 111 187 117
rect 191 111 195 117
rect 323 111 327 117
rect 331 111 335 117
rect 458 111 462 117
rect 466 111 470 117
rect 635 116 639 128
rect 653 116 657 128
rect 663 116 667 128
rect 681 116 685 128
rect 596 110 600 116
rect 604 110 608 116
rect 110 25 114 38
rect 128 25 132 38
rect 152 36 156 43
rect 160 36 164 43
rect 545 39 549 45
rect 553 39 557 45
rect 110 -49 114 -36
rect 128 -49 132 -36
rect 152 -38 156 -31
rect 160 -38 164 -31
rect 110 -118 114 -105
rect 128 -118 132 -105
rect 152 -107 156 -100
rect 160 -107 164 -100
rect 110 -192 114 -179
rect 128 -192 132 -179
rect 152 -181 156 -174
rect 160 -181 164 -174
rect 208 -229 212 31
rect 223 -229 228 31
rect 262 -228 266 32
rect 270 -228 274 32
rect 295 -228 299 32
rect 303 -228 307 32
rect 326 -228 330 32
rect 334 -228 338 32
rect 360 -227 364 33
rect 368 -227 372 33
rect 381 -227 385 33
rect 389 -227 393 33
rect 398 -227 402 33
rect 406 -227 410 33
rect 416 -226 420 34
rect 424 -226 428 34
rect 461 13 465 20
rect 469 13 473 20
rect 584 -10 588 2
rect 602 -10 606 2
rect 612 -10 616 2
rect 630 -10 634 2
rect 545 -16 549 -10
rect 553 -16 557 -10
rect 462 -72 466 -65
rect 470 -72 474 -65
rect 556 -97 560 -91
rect 564 -97 568 -91
rect 595 -146 599 -134
rect 613 -146 617 -134
rect 623 -146 627 -134
rect 641 -146 645 -134
rect 556 -152 560 -146
rect 564 -152 568 -146
rect 465 -183 469 -176
rect 473 -183 477 -176
rect 565 -231 569 -225
rect 573 -231 577 -225
rect 466 -255 470 -248
rect 474 -255 478 -248
rect 604 -280 608 -268
rect 622 -280 626 -268
rect 632 -280 636 -268
rect 650 -280 654 -268
rect 565 -286 569 -280
rect 573 -286 577 -280
rect 570 -380 574 -374
rect 578 -380 582 -374
rect 609 -429 613 -417
rect 627 -429 631 -417
rect 637 -429 641 -417
rect 655 -429 659 -417
rect 570 -435 574 -429
rect 578 -435 582 -429
<< pdcontact >>
rect 183 186 187 198
rect 191 186 195 198
rect 222 170 226 194
rect 231 170 235 194
rect 240 170 244 194
rect 250 164 254 188
rect 259 164 263 188
rect 268 164 272 188
rect 323 186 327 198
rect 331 186 335 198
rect 362 170 366 194
rect 371 170 375 194
rect 380 170 384 194
rect 183 131 187 143
rect 191 131 195 143
rect 390 164 394 188
rect 399 164 403 188
rect 408 164 412 188
rect 458 186 462 198
rect 466 186 470 198
rect 497 170 501 194
rect 506 170 510 194
rect 515 170 519 194
rect 323 131 327 143
rect 331 131 335 143
rect 525 164 529 188
rect 534 164 538 188
rect 543 164 547 188
rect 596 185 600 197
rect 604 185 608 197
rect 635 169 639 193
rect 644 169 648 193
rect 653 169 657 193
rect 458 131 462 143
rect 466 131 470 143
rect 663 163 667 187
rect 672 163 676 187
rect 681 163 685 187
rect 596 130 600 142
rect 604 130 608 142
rect 110 61 114 73
rect 119 61 123 73
rect 128 61 132 73
rect 152 61 156 73
rect 160 61 164 73
rect 215 63 219 75
rect 223 63 227 75
rect 251 63 255 75
rect 259 63 263 75
rect 292 63 296 75
rect 300 63 304 75
rect 327 63 331 75
rect 335 63 339 75
rect 545 59 549 71
rect 553 59 557 71
rect 461 38 465 50
rect 469 38 473 50
rect 584 43 588 67
rect 593 43 597 67
rect 602 43 606 67
rect 110 -13 114 -1
rect 119 -13 123 -1
rect 128 -13 132 -1
rect 152 -13 156 -1
rect 160 -13 164 -1
rect 110 -82 114 -70
rect 119 -82 123 -70
rect 128 -82 132 -70
rect 152 -82 156 -70
rect 160 -82 164 -70
rect 110 -156 114 -144
rect 119 -156 123 -144
rect 128 -156 132 -144
rect 152 -156 156 -144
rect 160 -156 164 -144
rect 612 37 616 61
rect 621 37 625 61
rect 630 37 634 61
rect 545 4 549 16
rect 553 4 557 16
rect 462 -47 466 -35
rect 470 -47 474 -35
rect 556 -77 560 -65
rect 564 -77 568 -65
rect 595 -93 599 -69
rect 604 -93 608 -69
rect 613 -93 617 -69
rect 623 -99 627 -75
rect 632 -99 636 -75
rect 641 -99 645 -75
rect 556 -132 560 -120
rect 564 -132 568 -120
rect 465 -158 469 -146
rect 473 -158 477 -146
rect 565 -211 569 -199
rect 573 -211 577 -199
rect 466 -230 470 -218
rect 474 -230 478 -218
rect 604 -227 608 -203
rect 613 -227 617 -203
rect 622 -227 626 -203
rect 632 -233 636 -209
rect 641 -233 645 -209
rect 650 -233 654 -209
rect 565 -266 569 -254
rect 573 -266 577 -254
rect 570 -360 574 -348
rect 578 -360 582 -348
rect 609 -376 613 -352
rect 618 -376 622 -352
rect 627 -376 631 -352
rect 637 -382 641 -358
rect 646 -382 650 -358
rect 655 -382 659 -358
rect 570 -415 574 -403
rect 578 -415 582 -403
<< polysilicon >>
rect 188 198 190 201
rect 328 198 330 201
rect 463 198 465 201
rect 227 194 229 197
rect 237 194 239 197
rect 188 172 190 186
rect 255 188 257 191
rect 265 188 267 191
rect 188 163 190 166
rect 227 161 229 170
rect 237 160 239 170
rect 367 194 369 197
rect 377 194 379 197
rect 328 172 330 186
rect 395 188 397 191
rect 405 188 407 191
rect 188 143 190 146
rect 188 117 190 131
rect 227 129 229 156
rect 237 129 239 155
rect 255 153 257 164
rect 255 129 257 149
rect 265 142 267 164
rect 328 163 330 166
rect 367 161 369 170
rect 377 160 379 170
rect 601 197 603 200
rect 502 194 504 197
rect 512 194 514 197
rect 463 172 465 186
rect 530 188 532 191
rect 540 188 542 191
rect 328 143 330 146
rect 265 129 267 138
rect 328 117 330 131
rect 367 129 369 156
rect 377 129 379 155
rect 395 153 397 164
rect 395 129 397 149
rect 405 142 407 164
rect 463 163 465 166
rect 502 161 504 170
rect 512 160 514 170
rect 640 193 642 196
rect 650 193 652 196
rect 601 171 603 185
rect 668 187 670 190
rect 678 187 680 190
rect 463 143 465 146
rect 405 129 407 138
rect 463 117 465 131
rect 502 129 504 156
rect 512 129 514 155
rect 530 153 532 164
rect 530 129 532 149
rect 540 142 542 164
rect 601 162 603 165
rect 640 160 642 169
rect 650 159 652 169
rect 601 142 603 145
rect 540 129 542 138
rect 227 114 229 117
rect 237 114 239 117
rect 255 114 257 117
rect 265 114 267 117
rect 367 114 369 117
rect 377 114 379 117
rect 395 114 397 117
rect 405 114 407 117
rect 502 114 504 117
rect 512 114 514 117
rect 530 114 532 117
rect 540 114 542 117
rect 601 116 603 130
rect 640 128 642 155
rect 650 128 652 154
rect 668 152 670 163
rect 668 128 670 148
rect 678 141 680 163
rect 678 128 680 137
rect 188 108 190 111
rect 328 108 330 111
rect 463 108 465 111
rect 640 113 642 116
rect 650 113 652 116
rect 668 113 670 116
rect 678 113 680 116
rect 601 107 603 110
rect 115 73 117 76
rect 125 73 127 76
rect 157 73 159 76
rect 220 75 222 78
rect 256 75 258 78
rect 297 75 299 78
rect 332 75 334 78
rect 550 71 552 74
rect 115 38 117 61
rect 125 38 127 61
rect 157 43 159 61
rect 220 48 222 63
rect 256 48 258 63
rect 297 48 299 63
rect 332 48 334 63
rect 589 67 591 70
rect 599 67 601 70
rect 466 50 468 53
rect 157 33 159 36
rect 213 31 215 39
rect 220 31 222 39
rect 267 32 269 39
rect 300 32 302 39
rect 331 32 333 39
rect 365 33 367 40
rect 386 33 388 40
rect 403 33 405 40
rect 421 34 423 41
rect 550 45 552 59
rect 617 61 619 64
rect 627 61 629 64
rect 115 21 117 25
rect 125 21 127 25
rect 115 -1 117 2
rect 125 -1 127 2
rect 157 -1 159 2
rect 115 -36 117 -13
rect 125 -36 127 -13
rect 157 -31 159 -13
rect 157 -41 159 -38
rect 115 -53 117 -49
rect 125 -53 127 -49
rect 115 -70 117 -67
rect 125 -70 127 -67
rect 157 -70 159 -67
rect 115 -105 117 -82
rect 125 -105 127 -82
rect 157 -100 159 -82
rect 157 -110 159 -107
rect 115 -122 117 -118
rect 125 -122 127 -118
rect 115 -144 117 -141
rect 125 -144 127 -141
rect 157 -144 159 -141
rect 115 -179 117 -156
rect 125 -179 127 -156
rect 157 -174 159 -156
rect 157 -184 159 -181
rect 115 -196 117 -192
rect 125 -196 127 -192
rect 466 20 468 38
rect 550 36 552 39
rect 589 34 591 43
rect 599 33 601 43
rect 550 16 552 19
rect 466 10 468 13
rect 550 -10 552 4
rect 589 2 591 29
rect 599 2 601 28
rect 617 26 619 37
rect 617 2 619 22
rect 627 15 629 37
rect 627 2 629 11
rect 589 -13 591 -10
rect 599 -13 601 -10
rect 617 -13 619 -10
rect 627 -13 629 -10
rect 550 -19 552 -16
rect 467 -35 469 -32
rect 467 -65 469 -47
rect 561 -65 563 -62
rect 467 -75 469 -72
rect 600 -69 602 -66
rect 610 -69 612 -66
rect 561 -91 563 -77
rect 628 -75 630 -72
rect 638 -75 640 -72
rect 561 -100 563 -97
rect 600 -102 602 -93
rect 610 -103 612 -93
rect 561 -120 563 -117
rect 470 -146 472 -143
rect 561 -146 563 -132
rect 600 -134 602 -107
rect 610 -134 612 -108
rect 628 -110 630 -99
rect 628 -134 630 -114
rect 638 -121 640 -99
rect 638 -134 640 -125
rect 600 -149 602 -146
rect 610 -149 612 -146
rect 628 -149 630 -146
rect 638 -149 640 -146
rect 561 -155 563 -152
rect 470 -176 472 -158
rect 470 -186 472 -183
rect 570 -199 572 -196
rect 609 -203 611 -200
rect 619 -203 621 -200
rect 471 -218 473 -215
rect 213 -232 215 -229
rect 220 -232 222 -229
rect 267 -232 269 -228
rect 300 -232 302 -228
rect 331 -232 333 -228
rect 365 -231 367 -227
rect 386 -231 388 -227
rect 403 -231 405 -227
rect 421 -230 423 -226
rect 570 -225 572 -211
rect 471 -248 473 -230
rect 637 -209 639 -206
rect 647 -209 649 -206
rect 570 -234 572 -231
rect 609 -236 611 -227
rect 619 -237 621 -227
rect 570 -254 572 -251
rect 471 -258 473 -255
rect 570 -280 572 -266
rect 609 -268 611 -241
rect 619 -268 621 -242
rect 637 -244 639 -233
rect 637 -268 639 -248
rect 647 -255 649 -233
rect 647 -268 649 -259
rect 609 -283 611 -280
rect 619 -283 621 -280
rect 637 -283 639 -280
rect 647 -283 649 -280
rect 570 -289 572 -286
rect 575 -348 577 -345
rect 614 -352 616 -349
rect 624 -352 626 -349
rect 575 -374 577 -360
rect 642 -358 644 -355
rect 652 -358 654 -355
rect 575 -383 577 -380
rect 614 -385 616 -376
rect 624 -386 626 -376
rect 575 -403 577 -400
rect 575 -429 577 -415
rect 614 -417 616 -390
rect 624 -417 626 -391
rect 642 -393 644 -382
rect 642 -417 644 -397
rect 652 -404 654 -382
rect 652 -417 654 -408
rect 614 -432 616 -429
rect 624 -432 626 -429
rect 642 -432 644 -429
rect 652 -432 654 -429
rect 575 -438 577 -435
<< polycontact >>
rect 184 175 188 179
rect 324 175 328 179
rect 184 120 188 124
rect 253 149 257 153
rect 459 175 463 179
rect 264 138 268 142
rect 324 120 328 124
rect 393 149 397 153
rect 597 174 601 178
rect 404 138 408 142
rect 459 120 463 124
rect 528 149 532 153
rect 539 138 543 142
rect 597 119 601 123
rect 666 148 670 152
rect 677 137 681 141
rect 111 48 115 52
rect 121 41 125 45
rect 153 47 157 51
rect 216 48 220 52
rect 252 48 256 52
rect 293 48 297 52
rect 328 48 332 52
rect 209 35 213 39
rect 222 35 226 39
rect 263 35 267 39
rect 296 35 300 39
rect 327 35 331 39
rect 361 36 365 40
rect 382 36 386 40
rect 399 36 403 40
rect 417 37 421 41
rect 546 48 550 52
rect 111 -26 115 -22
rect 121 -33 125 -29
rect 153 -27 157 -23
rect 111 -95 115 -91
rect 121 -102 125 -98
rect 153 -96 157 -92
rect 111 -169 115 -165
rect 121 -176 125 -172
rect 153 -170 157 -166
rect 462 24 466 28
rect 546 -7 550 -3
rect 615 22 619 26
rect 626 11 630 15
rect 463 -61 467 -57
rect 557 -88 561 -84
rect 557 -143 561 -139
rect 626 -114 630 -110
rect 637 -125 641 -121
rect 466 -172 470 -168
rect 566 -222 570 -218
rect 467 -244 471 -240
rect 566 -277 570 -273
rect 635 -248 639 -244
rect 646 -259 650 -255
rect 571 -371 575 -367
rect 571 -426 575 -422
rect 640 -397 644 -393
rect 651 -408 655 -404
<< metal1 >>
rect 182 204 210 207
rect 322 204 350 207
rect 457 204 485 207
rect 183 198 186 204
rect 207 203 210 204
rect 207 200 278 203
rect 166 174 169 177
rect 174 175 184 178
rect 192 178 195 186
rect 222 194 225 200
rect 241 194 244 200
rect 323 198 326 204
rect 347 203 350 204
rect 347 200 418 203
rect 192 175 213 178
rect 192 172 195 175
rect 183 162 186 166
rect 177 160 201 162
rect 177 159 195 160
rect 200 159 201 160
rect 210 152 213 175
rect 251 194 271 197
rect 251 188 254 194
rect 268 188 271 194
rect 232 167 235 170
rect 232 164 250 167
rect 306 174 309 177
rect 314 175 324 178
rect 332 178 335 186
rect 362 194 365 200
rect 381 194 384 200
rect 458 198 461 204
rect 482 203 485 204
rect 595 203 623 206
rect 482 200 553 203
rect 332 175 353 178
rect 332 172 335 175
rect 260 157 263 164
rect 323 162 326 166
rect 317 160 341 162
rect 317 159 335 160
rect 260 154 277 157
rect 182 151 201 152
rect 177 149 201 151
rect 210 149 253 152
rect 183 143 186 149
rect 274 143 277 154
rect 340 159 341 160
rect 350 152 353 175
rect 391 194 411 197
rect 391 188 394 194
rect 408 188 411 194
rect 372 167 375 170
rect 372 164 390 167
rect 441 174 444 177
rect 449 175 459 178
rect 467 178 470 186
rect 497 194 500 200
rect 516 194 519 200
rect 596 197 599 203
rect 620 202 623 203
rect 620 199 691 202
rect 467 175 488 178
rect 467 172 470 175
rect 400 157 403 164
rect 458 162 461 166
rect 452 160 476 162
rect 452 159 470 160
rect 400 154 417 157
rect 322 151 341 152
rect 317 149 341 151
rect 350 149 393 152
rect 323 143 326 149
rect 414 143 417 154
rect 475 159 476 160
rect 485 152 488 175
rect 526 194 546 197
rect 526 188 529 194
rect 543 188 546 194
rect 507 167 510 170
rect 507 164 525 167
rect 579 173 582 176
rect 587 174 597 177
rect 605 177 608 185
rect 635 193 638 199
rect 654 193 657 199
rect 605 174 626 177
rect 605 171 608 174
rect 535 157 538 164
rect 596 161 599 165
rect 590 159 614 161
rect 590 158 608 159
rect 535 154 552 157
rect 457 151 476 152
rect 452 149 476 151
rect 485 149 528 152
rect 458 143 461 149
rect 549 143 552 154
rect 613 158 614 159
rect 623 151 626 174
rect 664 193 684 196
rect 664 187 667 193
rect 681 187 684 193
rect 645 166 648 169
rect 645 163 663 166
rect 673 156 676 163
rect 673 153 690 156
rect 595 150 614 151
rect 590 148 614 150
rect 623 148 666 151
rect 239 138 264 141
rect 274 139 287 143
rect 239 136 242 138
rect 166 120 169 123
rect 174 120 184 123
rect 192 123 195 131
rect 204 133 242 136
rect 274 135 277 139
rect 204 123 207 133
rect 245 132 277 135
rect 245 129 248 132
rect 192 120 207 123
rect 192 117 195 120
rect 244 126 250 129
rect 183 107 186 111
rect 204 110 209 113
rect 222 113 225 117
rect 269 113 272 117
rect 214 110 278 113
rect 204 107 207 110
rect 177 104 207 107
rect 283 99 287 139
rect 379 138 404 141
rect 414 139 426 143
rect 379 136 382 138
rect 306 120 309 123
rect 314 120 324 123
rect 332 123 335 131
rect 344 133 382 136
rect 414 135 417 139
rect 344 123 347 133
rect 385 132 417 135
rect 385 129 388 132
rect 332 120 347 123
rect 332 117 335 120
rect 384 126 390 129
rect 323 107 326 111
rect 344 110 349 113
rect 362 113 365 117
rect 409 113 412 117
rect 354 110 418 113
rect 344 107 347 110
rect 317 104 347 107
rect 422 98 426 139
rect 514 138 539 141
rect 549 139 560 143
rect 514 136 517 138
rect 441 120 444 123
rect 449 120 459 123
rect 467 123 470 131
rect 479 133 517 136
rect 549 135 552 139
rect 479 123 482 133
rect 520 132 552 135
rect 520 129 523 132
rect 467 120 482 123
rect 467 117 470 120
rect 519 126 525 129
rect 458 107 461 111
rect 479 110 484 113
rect 497 113 500 117
rect 544 113 547 117
rect 489 110 553 113
rect 479 107 482 110
rect 452 104 482 107
rect 556 99 560 139
rect 596 142 599 148
rect 687 142 690 153
rect 652 137 677 140
rect 687 138 702 142
rect 652 135 655 137
rect 579 119 582 122
rect 587 119 597 122
rect 605 122 608 130
rect 617 132 655 135
rect 687 134 690 138
rect 617 122 620 132
rect 658 131 690 134
rect 658 128 661 131
rect 605 119 620 122
rect 605 116 608 119
rect 657 125 663 128
rect 596 106 599 110
rect 617 109 622 112
rect 635 112 638 116
rect 682 112 685 116
rect 627 109 691 112
rect 617 106 620 109
rect 590 103 620 106
rect 698 100 702 138
rect 422 94 429 98
rect 553 95 560 99
rect 102 79 173 82
rect 208 81 236 84
rect 244 81 272 84
rect 285 81 313 84
rect 320 81 348 84
rect 110 73 114 79
rect 128 73 132 79
rect 152 73 155 79
rect 215 75 218 81
rect 251 75 254 81
rect 292 75 295 81
rect 327 75 330 81
rect 544 77 572 80
rect 119 58 122 61
rect 119 55 132 58
rect 102 48 111 52
rect 129 51 132 55
rect 161 51 164 61
rect 129 47 153 51
rect 161 48 173 51
rect 208 48 216 52
rect 224 48 227 63
rect 244 48 252 52
rect 260 48 263 63
rect 285 48 293 52
rect 301 48 304 63
rect 320 48 328 52
rect 336 48 339 63
rect 545 71 548 77
rect 569 76 572 77
rect 569 73 640 76
rect 450 56 482 59
rect 461 50 464 56
rect 102 41 121 45
rect 129 38 132 47
rect 161 43 164 48
rect 110 19 113 25
rect 152 19 155 36
rect 206 35 209 39
rect 226 35 232 39
rect 260 35 263 39
rect 293 35 296 39
rect 324 35 327 39
rect 334 32 338 39
rect 358 36 361 40
rect 368 33 372 40
rect 379 36 382 40
rect 389 33 393 40
rect 396 36 399 40
rect 406 33 410 40
rect 414 37 417 41
rect 424 34 428 41
rect 528 47 531 50
rect 536 48 546 51
rect 554 51 557 59
rect 584 67 587 73
rect 603 67 606 73
rect 554 48 575 51
rect 554 45 557 48
rect 102 16 155 19
rect 102 5 173 8
rect 110 -1 114 5
rect 128 -1 132 5
rect 152 -1 155 5
rect 119 -16 122 -13
rect 119 -19 132 -16
rect 102 -26 111 -22
rect 129 -23 132 -19
rect 161 -23 164 -13
rect 129 -27 153 -23
rect 161 -26 173 -23
rect 102 -33 121 -29
rect 129 -36 132 -27
rect 161 -31 164 -26
rect 110 -55 113 -49
rect 152 -55 155 -38
rect 102 -58 155 -55
rect 102 -64 173 -61
rect 110 -70 114 -64
rect 128 -70 132 -64
rect 152 -70 155 -64
rect 119 -85 122 -82
rect 119 -88 132 -85
rect 102 -95 111 -91
rect 129 -92 132 -88
rect 161 -92 164 -82
rect 129 -96 153 -92
rect 161 -95 173 -92
rect 102 -102 121 -98
rect 129 -105 132 -96
rect 161 -100 164 -95
rect 110 -124 113 -118
rect 152 -124 155 -107
rect 102 -127 155 -124
rect 102 -138 173 -135
rect 110 -144 114 -138
rect 128 -144 132 -138
rect 152 -144 155 -138
rect 119 -159 122 -156
rect 119 -162 132 -159
rect 102 -169 111 -165
rect 129 -166 132 -162
rect 161 -166 164 -156
rect 129 -170 153 -166
rect 161 -169 173 -166
rect 102 -176 121 -172
rect 129 -179 132 -170
rect 161 -174 164 -169
rect 110 -198 113 -192
rect 152 -198 155 -181
rect 102 -201 155 -198
rect 208 -238 212 -229
rect 223 -230 228 -229
rect 262 -230 266 -228
rect 223 -235 266 -230
rect 270 -230 274 -228
rect 295 -230 299 -228
rect 270 -235 299 -230
rect 303 -230 307 -228
rect 470 28 473 38
rect 545 35 548 39
rect 539 33 563 35
rect 539 32 557 33
rect 450 24 462 28
rect 470 25 482 28
rect 470 20 473 25
rect 562 32 563 33
rect 572 25 575 48
rect 613 67 633 70
rect 613 61 616 67
rect 630 61 633 67
rect 594 40 597 43
rect 594 37 612 40
rect 622 30 625 37
rect 622 27 639 30
rect 544 24 563 25
rect 539 22 563 24
rect 572 22 615 25
rect 545 16 548 22
rect 636 16 639 27
rect 461 -4 464 13
rect 601 11 626 14
rect 636 12 649 16
rect 601 9 604 11
rect 450 -7 464 -4
rect 528 -7 531 -4
rect 536 -7 546 -4
rect 554 -4 557 4
rect 566 6 604 9
rect 636 8 639 12
rect 566 -4 569 6
rect 607 5 639 8
rect 607 2 610 5
rect 554 -7 569 -4
rect 554 -10 557 -7
rect 606 -1 612 2
rect 545 -20 548 -16
rect 566 -17 571 -14
rect 584 -14 587 -10
rect 631 -14 634 -10
rect 576 -17 640 -14
rect 566 -20 569 -17
rect 539 -23 569 -20
rect 451 -29 483 -26
rect 645 -28 649 12
rect 462 -35 465 -29
rect 471 -57 474 -47
rect 451 -61 463 -57
rect 471 -60 483 -57
rect 555 -59 583 -56
rect 471 -65 474 -60
rect 556 -65 559 -59
rect 580 -60 583 -59
rect 580 -63 651 -60
rect 462 -89 465 -72
rect 539 -89 542 -86
rect 451 -92 465 -89
rect 547 -88 557 -85
rect 565 -85 568 -77
rect 595 -69 598 -63
rect 614 -69 617 -63
rect 565 -88 586 -85
rect 565 -91 568 -88
rect 556 -101 559 -97
rect 550 -103 574 -101
rect 550 -104 568 -103
rect 573 -104 574 -103
rect 583 -111 586 -88
rect 624 -69 644 -66
rect 624 -75 627 -69
rect 641 -75 644 -69
rect 605 -96 608 -93
rect 605 -99 623 -96
rect 633 -106 636 -99
rect 633 -109 650 -106
rect 555 -112 574 -111
rect 550 -114 574 -112
rect 583 -114 626 -111
rect 556 -120 559 -114
rect 647 -120 650 -109
rect 612 -125 637 -122
rect 647 -124 660 -120
rect 612 -127 615 -125
rect 454 -140 486 -137
rect 465 -146 468 -140
rect 539 -143 542 -140
rect 547 -143 557 -140
rect 565 -140 568 -132
rect 577 -130 615 -127
rect 647 -128 650 -124
rect 577 -140 580 -130
rect 618 -131 650 -128
rect 618 -134 621 -131
rect 565 -143 580 -140
rect 565 -146 568 -143
rect 617 -137 623 -134
rect 556 -156 559 -152
rect 577 -153 582 -150
rect 595 -150 598 -146
rect 642 -150 645 -146
rect 587 -153 651 -150
rect 577 -156 580 -153
rect 474 -168 477 -158
rect 550 -159 580 -156
rect 656 -164 660 -124
rect 454 -172 466 -168
rect 474 -171 486 -168
rect 474 -176 477 -171
rect 465 -200 468 -183
rect 564 -193 592 -190
rect 454 -203 468 -200
rect 565 -199 568 -193
rect 589 -194 592 -193
rect 589 -197 660 -194
rect 455 -212 487 -209
rect 466 -218 469 -212
rect 326 -230 330 -228
rect 303 -235 330 -230
rect 360 -232 364 -227
rect 381 -232 385 -227
rect 398 -232 402 -227
rect 416 -232 420 -226
rect 548 -223 551 -220
rect 556 -222 566 -219
rect 574 -219 577 -211
rect 604 -203 607 -197
rect 623 -203 626 -197
rect 574 -222 595 -219
rect 574 -225 577 -222
rect 360 -235 420 -232
rect 203 -242 221 -238
rect 475 -240 478 -230
rect 565 -235 568 -231
rect 559 -237 583 -235
rect 559 -238 577 -237
rect 455 -244 467 -240
rect 475 -243 487 -240
rect 475 -248 478 -243
rect 582 -238 583 -237
rect 592 -245 595 -222
rect 633 -203 653 -200
rect 633 -209 636 -203
rect 650 -209 653 -203
rect 614 -230 617 -227
rect 614 -233 632 -230
rect 642 -240 645 -233
rect 642 -243 659 -240
rect 564 -246 583 -245
rect 559 -248 583 -246
rect 592 -248 635 -245
rect 565 -254 568 -248
rect 656 -254 659 -243
rect 466 -272 469 -255
rect 621 -259 646 -256
rect 656 -258 669 -254
rect 621 -261 624 -259
rect 455 -275 469 -272
rect 548 -277 551 -274
rect 556 -277 566 -274
rect 574 -274 577 -266
rect 586 -264 624 -261
rect 656 -262 659 -258
rect 586 -274 589 -264
rect 627 -265 659 -262
rect 627 -268 630 -265
rect 574 -277 589 -274
rect 574 -280 577 -277
rect 626 -271 632 -268
rect 565 -290 568 -286
rect 586 -287 591 -284
rect 604 -284 607 -280
rect 651 -284 654 -280
rect 596 -287 660 -284
rect 586 -290 589 -287
rect 559 -293 589 -290
rect 665 -298 669 -258
rect 569 -342 597 -339
rect 570 -348 573 -342
rect 594 -343 597 -342
rect 594 -346 665 -343
rect 553 -372 556 -369
rect 561 -371 571 -368
rect 579 -368 582 -360
rect 609 -352 612 -346
rect 628 -352 631 -346
rect 579 -371 600 -368
rect 579 -374 582 -371
rect 570 -384 573 -380
rect 564 -386 588 -384
rect 564 -387 582 -386
rect 587 -387 588 -386
rect 597 -394 600 -371
rect 638 -352 658 -349
rect 638 -358 641 -352
rect 655 -358 658 -352
rect 619 -379 622 -376
rect 619 -382 637 -379
rect 647 -389 650 -382
rect 647 -392 664 -389
rect 569 -395 588 -394
rect 564 -397 588 -395
rect 597 -397 640 -394
rect 570 -403 573 -397
rect 661 -403 664 -392
rect 626 -408 651 -405
rect 661 -407 674 -403
rect 626 -410 629 -408
rect 553 -426 556 -423
rect 561 -426 571 -423
rect 579 -423 582 -415
rect 591 -413 629 -410
rect 661 -411 664 -407
rect 591 -423 594 -413
rect 632 -414 664 -411
rect 632 -417 635 -414
rect 579 -426 594 -423
rect 579 -429 582 -426
rect 631 -420 637 -417
rect 570 -439 573 -435
rect 591 -436 596 -433
rect 609 -433 612 -429
rect 656 -433 659 -429
rect 601 -436 665 -433
rect 591 -439 594 -436
rect 564 -442 594 -439
rect 670 -447 674 -407
<< m2contact >>
rect 169 173 174 178
rect 309 173 314 178
rect 444 173 449 178
rect 582 172 587 177
rect 169 119 174 124
rect 309 119 314 124
rect 444 119 449 124
rect 582 118 587 123
rect 531 46 536 51
rect 531 -8 536 -3
rect 542 -90 547 -85
rect 542 -144 547 -139
rect 551 -224 556 -219
rect 551 -278 556 -273
rect 556 -373 561 -368
rect 556 -427 561 -422
<< pm12contact >>
rect 225 156 230 161
rect 234 155 239 160
rect 365 156 370 161
rect 374 155 379 160
rect 500 156 505 161
rect 509 155 514 160
rect 638 155 643 160
rect 647 154 652 159
rect 587 29 592 34
rect 596 28 601 33
rect 598 -107 603 -102
rect 607 -108 612 -103
rect 607 -241 612 -236
rect 616 -242 621 -237
rect 612 -390 617 -385
rect 621 -391 626 -386
<< metal2 >>
rect 170 167 173 173
rect 310 167 313 173
rect 445 167 448 173
rect 170 164 207 167
rect 310 164 347 167
rect 445 164 482 167
rect 204 161 207 164
rect 344 161 347 164
rect 479 161 482 164
rect 583 166 586 172
rect 583 163 620 166
rect 204 158 225 161
rect 234 145 237 155
rect 344 158 365 161
rect 374 145 377 155
rect 479 158 500 161
rect 617 160 620 163
rect 509 145 512 155
rect 617 157 638 160
rect 171 142 237 145
rect 311 142 377 145
rect 446 142 512 145
rect 647 144 650 154
rect 171 124 174 142
rect 311 124 314 142
rect 446 124 449 142
rect 584 141 650 144
rect 584 123 587 141
rect 532 40 535 46
rect 532 37 569 40
rect 566 34 569 37
rect 566 31 587 34
rect 596 18 599 28
rect 533 15 599 18
rect 533 -3 536 15
rect 543 -96 546 -90
rect 543 -99 580 -96
rect 577 -102 580 -99
rect 577 -105 598 -102
rect 607 -118 610 -108
rect 544 -121 610 -118
rect 544 -139 547 -121
rect 552 -230 555 -224
rect 552 -233 589 -230
rect 586 -236 589 -233
rect 586 -239 607 -236
rect 616 -252 619 -242
rect 553 -255 619 -252
rect 553 -273 556 -255
rect 557 -379 560 -373
rect 557 -382 594 -379
rect 591 -385 594 -382
rect 591 -388 612 -385
rect 621 -401 624 -391
rect 558 -404 624 -401
rect 558 -422 561 -404
<< m123contact >>
rect 177 204 182 209
rect 317 204 322 209
rect 452 204 457 209
rect 590 203 595 208
rect 177 151 182 156
rect 195 155 200 160
rect 317 151 322 156
rect 335 155 340 160
rect 452 151 457 156
rect 470 155 475 160
rect 590 150 595 155
rect 608 154 613 159
rect 209 110 214 115
rect 349 110 354 115
rect 484 110 489 115
rect 622 109 627 114
rect 539 77 544 82
rect 539 24 544 29
rect 557 28 562 33
rect 571 -17 576 -12
rect 550 -59 555 -54
rect 550 -112 555 -107
rect 568 -108 573 -103
rect 582 -153 587 -148
rect 559 -193 564 -188
rect 559 -246 564 -241
rect 577 -242 582 -237
rect 591 -287 596 -282
rect 564 -342 569 -337
rect 564 -395 569 -390
rect 582 -391 587 -386
rect 596 -436 601 -431
<< metal3 >>
rect 177 156 180 204
rect 200 155 212 158
rect 209 115 212 155
rect 317 156 320 204
rect 340 155 352 158
rect 349 115 352 155
rect 452 156 455 204
rect 475 155 487 158
rect 484 115 487 155
rect 590 155 593 203
rect 613 154 625 157
rect 622 114 625 154
rect 539 29 542 77
rect 562 28 574 31
rect 571 -12 574 28
rect 550 -107 553 -59
rect 573 -108 585 -105
rect 582 -148 585 -108
rect 559 -241 562 -193
rect 582 -242 594 -239
rect 591 -282 594 -242
rect 564 -390 567 -342
rect 587 -391 599 -388
rect 596 -431 599 -391
<< labels >>
rlabel metal1 195 104 199 107 1 gnd
rlabel metal1 245 110 248 112 1 gnd
rlabel metal1 193 160 194 162 1 gnd
rlabel metal1 189 204 192 206 5 vdd
rlabel metal1 190 150 193 152 1 vdd
rlabel metal1 274 139 278 143 7 p0
rlabel metal1 166 174 167 177 1 a0
rlabel metal1 166 120 167 123 1 b0
rlabel metal1 335 104 339 107 1 gnd
rlabel metal1 385 110 388 112 1 gnd
rlabel metal1 333 160 334 162 1 gnd
rlabel metal1 329 204 332 206 5 vdd
rlabel metal1 330 150 333 152 1 vdd
rlabel metal1 470 104 474 107 1 gnd
rlabel metal1 520 110 523 112 1 gnd
rlabel metal1 468 160 469 162 1 gnd
rlabel metal1 464 204 467 206 5 vdd
rlabel metal1 465 150 468 152 1 vdd
rlabel metal1 608 103 612 106 1 gnd
rlabel metal1 658 109 661 111 1 gnd
rlabel metal1 606 159 607 161 1 gnd
rlabel metal1 602 203 605 205 5 vdd
rlabel metal1 603 149 606 151 1 vdd
rlabel metal1 306 120 307 123 1 b1
rlabel metal1 306 174 307 177 1 a1
rlabel metal1 441 174 442 177 1 a2
rlabel metal1 441 120 442 123 1 b2
rlabel metal1 579 173 580 176 1 a3
rlabel metal1 579 119 580 122 1 b3
rlabel metal1 687 138 691 142 7 p3
rlabel metal1 414 139 418 143 1 p1
rlabel metal1 549 139 553 143 1 p2
rlabel metal1 168 49 169 50 7 g0
rlabel metal1 105 43 106 44 3 b0
rlabel metal1 103 50 104 51 3 a0
rlabel metal1 128 17 128 17 1 gnd!
rlabel metal1 128 81 128 81 5 vdd!
rlabel metal1 168 -25 169 -24 7 g1
rlabel metal1 128 -126 128 -126 1 gnd!
rlabel metal1 128 -62 128 -62 5 vdd!
rlabel metal1 128 -200 128 -200 1 gnd!
rlabel metal1 128 -136 128 -136 5 vdd!
rlabel metal1 103 -93 104 -92 3 a2
rlabel metal1 105 -100 106 -99 3 b2
rlabel metal1 104 -167 105 -166 3 a3
rlabel metal1 105 -174 106 -173 3 b3
rlabel metal1 168 -168 169 -167 7 g3
rlabel metal1 105 -31 106 -30 3 b1
rlabel metal1 104 -24 105 -23 3 a1
rlabel metal1 128 7 128 7 5 vdd!
rlabel metal1 128 -57 128 -57 1 gnd!
rlabel metal1 221 82 228 83 1 vdd
rlabel metal1 210 49 213 51 1 gnd
rlabel metal1 225 50 226 51 1 c3b
rlabel metal1 207 36 208 37 1 cin
rlabel metal1 228 36 229 38 1 p0
rlabel metal1 257 82 264 83 1 vdd
rlabel metal1 246 49 249 51 1 gnd
rlabel metal1 298 82 305 83 1 vdd
rlabel metal1 287 49 290 51 1 gnd
rlabel metal1 333 82 340 83 1 vdd
rlabel metal1 322 49 325 51 1 gnd
rlabel metal1 261 50 262 51 1 c2b
rlabel metal1 302 50 303 51 1 c1b
rlabel metal1 337 50 338 51 1 c0b
rlabel metal1 261 36 262 37 1 p1
rlabel metal1 294 36 295 37 1 p2
rlabel metal1 325 36 326 37 1 p3
rlabel metal1 335 35 337 37 1 c3b
rlabel metal1 359 37 360 38 1 g0
rlabel metal1 369 36 371 38 1 c0b
rlabel metal1 380 37 381 38 1 g1
rlabel metal1 390 36 392 38 1 c1b
rlabel metal1 397 37 398 38 1 g2
rlabel metal1 407 36 409 38 1 c2b
rlabel metal1 415 38 416 39 1 g3
rlabel metal1 425 37 427 39 1 c3b
rlabel metal1 557 -23 561 -20 1 gnd
rlabel metal1 607 -17 610 -15 1 gnd
rlabel metal1 555 33 556 35 1 gnd
rlabel metal1 551 77 554 79 5 vdd
rlabel metal1 552 23 555 25 1 vdd
rlabel metal1 568 -159 572 -156 1 gnd
rlabel metal1 618 -153 621 -151 1 gnd
rlabel metal1 566 -103 567 -101 1 gnd
rlabel metal1 562 -59 565 -57 5 vdd
rlabel metal1 563 -113 566 -111 1 vdd
rlabel metal1 577 -293 581 -290 1 gnd
rlabel metal1 627 -287 630 -285 1 gnd
rlabel metal1 575 -237 576 -235 1 gnd
rlabel metal1 571 -193 574 -191 5 vdd
rlabel metal1 572 -247 575 -245 1 vdd
rlabel metal1 582 -442 586 -439 1 gnd
rlabel metal1 632 -436 635 -434 1 gnd
rlabel metal1 580 -386 581 -384 1 gnd
rlabel metal1 576 -342 579 -340 5 vdd
rlabel metal1 577 -396 580 -394 1 vdd
rlabel metal1 528 47 529 50 1 p0
rlabel metal1 528 -7 529 -4 1 cin
rlabel metal1 636 12 640 16 1 s0
rlabel metal1 539 -89 540 -86 1 p1
rlabel metal1 539 -143 540 -140 1 c0
rlabel metal1 647 -124 651 -120 1 s1
rlabel metal1 548 -223 549 -220 1 p2
rlabel metal1 548 -277 549 -274 1 c1
rlabel metal1 656 -258 660 -254 1 s2
rlabel metal1 553 -372 554 -369 1 p3
rlabel metal1 553 -426 554 -423 1 c2
rlabel metal1 661 -407 665 -403 1 s3
rlabel metal1 168 -94 169 -93 7 g2
rlabel metal1 453 25 454 27 1 c0b
rlabel metal1 455 -60 458 -58 1 c1b
rlabel metal1 459 -171 462 -169 1 c2b
rlabel metal1 460 -243 463 -241 1 c3b
rlabel metal1 477 26 480 28 1 c0
rlabel metal1 478 -59 479 -58 1 c1
rlabel metal1 481 -170 482 -169 1 c2
rlabel metal1 482 -242 483 -241 1 c3
rlabel metal1 460 -274 462 -273 1 gnd
rlabel metal1 467 -211 469 -210 1 vdd
rlabel metal1 460 -201 462 -200 1 gnd
rlabel metal1 466 -139 468 -138 1 vdd
rlabel metal1 457 -91 459 -90 1 gnd
rlabel metal1 465 -28 467 -27 1 vdd
rlabel metal1 454 -6 456 -5 1 gnd
rlabel metal1 462 57 464 58 1 vdd
rlabel metal1 212 -241 218 -239 1 gnd
rlabel metal1 240 -235 247 -230 1 c0b
rlabel metal1 279 -235 286 -230 1 c1b
rlabel metal1 314 -235 321 -230 1 c2b
rlabel metal1 383 -235 386 -233 1 gnd
<< end >>
